VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO tristate_inv_delay_line_128
  CLASS BLOCK ;
  ORIGIN 2.88 3 ;
  FOREIGN tristate_inv_delay_line_128 -2.88 -3 ;
  SIZE 772.825 BY 12.92 ;
  SYMMETRY X Y R90 ;
  PIN clk_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT -1.47 9.6 -1.15 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT -1.47 -3 -1.15 -2.68 ;
    END
  END clk_in
  PIN clk_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.52 9.6 1.84 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.52 -3 1.84 -2.68 ;
    END
  END clk_out
  PIN ctl[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.03 9.6 0.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.03 -3 0.35 -2.68 ;
    END
  END ctl[0]
  PIN ctl[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 600.03 9.6 600.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 600.03 -3 600.35 -2.68 ;
    END
  END ctl[100]
  PIN ctl[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 606.03 9.6 606.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 606.03 -3 606.35 -2.68 ;
    END
  END ctl[101]
  PIN ctl[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 612.03 9.6 612.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 612.03 -3 612.35 -2.68 ;
    END
  END ctl[102]
  PIN ctl[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 618.03 9.6 618.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 618.03 -3 618.35 -2.68 ;
    END
  END ctl[103]
  PIN ctl[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 624.03 9.6 624.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 624.03 -3 624.35 -2.68 ;
    END
  END ctl[104]
  PIN ctl[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 630.03 9.6 630.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 630.03 -3 630.35 -2.68 ;
    END
  END ctl[105]
  PIN ctl[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 636.03 9.6 636.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 636.03 -3 636.35 -2.68 ;
    END
  END ctl[106]
  PIN ctl[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 642.03 9.6 642.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 642.03 -3 642.35 -2.68 ;
    END
  END ctl[107]
  PIN ctl[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 648.03 9.6 648.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 648.03 -3 648.35 -2.68 ;
    END
  END ctl[108]
  PIN ctl[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 654.03 9.6 654.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 654.03 -3 654.35 -2.68 ;
    END
  END ctl[109]
  PIN ctl[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 60.03 9.6 60.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 60.03 -3 60.35 -2.68 ;
    END
  END ctl[10]
  PIN ctl[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 660.03 9.6 660.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 660.03 -3 660.35 -2.68 ;
    END
  END ctl[110]
  PIN ctl[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 666.03 9.6 666.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 666.03 -3 666.35 -2.68 ;
    END
  END ctl[111]
  PIN ctl[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 672.03 9.6 672.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 672.03 -3 672.35 -2.68 ;
    END
  END ctl[112]
  PIN ctl[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 678.03 9.6 678.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 678.03 -3 678.35 -2.68 ;
    END
  END ctl[113]
  PIN ctl[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 684.03 9.6 684.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 684.03 -3 684.35 -2.68 ;
    END
  END ctl[114]
  PIN ctl[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 690.03 9.6 690.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 690.03 -3 690.35 -2.68 ;
    END
  END ctl[115]
  PIN ctl[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 696.03 9.6 696.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 696.03 -3 696.35 -2.68 ;
    END
  END ctl[116]
  PIN ctl[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 702.03 9.6 702.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 702.03 -3 702.35 -2.68 ;
    END
  END ctl[117]
  PIN ctl[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 708.03 9.6 708.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 708.03 -3 708.35 -2.68 ;
    END
  END ctl[118]
  PIN ctl[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 714.03 9.6 714.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 714.03 -3 714.35 -2.68 ;
    END
  END ctl[119]
  PIN ctl[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 66.03 9.6 66.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 66.03 -3 66.35 -2.68 ;
    END
  END ctl[11]
  PIN ctl[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 720.03 9.6 720.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 720.03 -3 720.35 -2.68 ;
    END
  END ctl[120]
  PIN ctl[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 726.03 9.6 726.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 726.03 -3 726.35 -2.68 ;
    END
  END ctl[121]
  PIN ctl[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 732.03 9.6 732.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 732.03 -3 732.35 -2.68 ;
    END
  END ctl[122]
  PIN ctl[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 738.03 9.6 738.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 738.03 -3 738.35 -2.68 ;
    END
  END ctl[123]
  PIN ctl[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 744.03 9.6 744.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 744.03 -3 744.35 -2.68 ;
    END
  END ctl[124]
  PIN ctl[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 750.03 9.6 750.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 750.03 -3 750.35 -2.68 ;
    END
  END ctl[125]
  PIN ctl[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 756.03 9.6 756.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 756.03 -3 756.35 -2.68 ;
    END
  END ctl[126]
  PIN ctl[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 762.03 9.6 762.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 762.03 -3 762.35 -2.68 ;
    END
  END ctl[127]
  PIN ctl[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 72.03 9.6 72.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 72.03 -3 72.35 -2.68 ;
    END
  END ctl[12]
  PIN ctl[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 78.03 9.6 78.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 78.03 -3 78.35 -2.68 ;
    END
  END ctl[13]
  PIN ctl[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 84.03 9.6 84.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 84.03 -3 84.35 -2.68 ;
    END
  END ctl[14]
  PIN ctl[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 90.03 9.6 90.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 90.03 -3 90.35 -2.68 ;
    END
  END ctl[15]
  PIN ctl[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 96.03 9.6 96.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 96.03 -3 96.35 -2.68 ;
    END
  END ctl[16]
  PIN ctl[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 102.03 9.6 102.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 102.03 -3 102.35 -2.68 ;
    END
  END ctl[17]
  PIN ctl[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 108.03 9.6 108.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 108.03 -3 108.35 -2.68 ;
    END
  END ctl[18]
  PIN ctl[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 114.03 9.6 114.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 114.03 -3 114.35 -2.68 ;
    END
  END ctl[19]
  PIN ctl[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 6.03 9.6 6.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.03 -3 6.35 -2.68 ;
    END
  END ctl[1]
  PIN ctl[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 120.03 9.6 120.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 120.03 -3 120.35 -2.68 ;
    END
  END ctl[20]
  PIN ctl[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 126.03 9.6 126.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 126.03 -3 126.35 -2.68 ;
    END
  END ctl[21]
  PIN ctl[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 132.03 9.6 132.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 132.03 -3 132.35 -2.68 ;
    END
  END ctl[22]
  PIN ctl[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 138.03 9.6 138.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 138.03 -3 138.35 -2.68 ;
    END
  END ctl[23]
  PIN ctl[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 144.03 9.6 144.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 144.03 -3 144.35 -2.68 ;
    END
  END ctl[24]
  PIN ctl[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 150.03 9.6 150.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 150.03 -3 150.35 -2.68 ;
    END
  END ctl[25]
  PIN ctl[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 156.03 9.6 156.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 156.03 -3 156.35 -2.68 ;
    END
  END ctl[26]
  PIN ctl[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 162.03 9.6 162.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 162.03 -3 162.35 -2.68 ;
    END
  END ctl[27]
  PIN ctl[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 168.03 9.6 168.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 168.03 -3 168.35 -2.68 ;
    END
  END ctl[28]
  PIN ctl[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 174.03 9.6 174.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 174.03 -3 174.35 -2.68 ;
    END
  END ctl[29]
  PIN ctl[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 12.03 9.6 12.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 12.03 -3 12.35 -2.68 ;
    END
  END ctl[2]
  PIN ctl[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 180.03 9.6 180.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 180.03 -3 180.35 -2.68 ;
    END
  END ctl[30]
  PIN ctl[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 186.03 9.6 186.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 186.03 -3 186.35 -2.68 ;
    END
  END ctl[31]
  PIN ctl[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 192.03 9.6 192.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 192.03 -3 192.35 -2.68 ;
    END
  END ctl[32]
  PIN ctl[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 198.03 9.6 198.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 198.03 -3 198.35 -2.68 ;
    END
  END ctl[33]
  PIN ctl[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 204.03 9.6 204.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 204.03 -3 204.35 -2.68 ;
    END
  END ctl[34]
  PIN ctl[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 210.03 9.6 210.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 210.03 -3 210.35 -2.68 ;
    END
  END ctl[35]
  PIN ctl[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 216.03 9.6 216.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 216.03 -3 216.35 -2.68 ;
    END
  END ctl[36]
  PIN ctl[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 222.03 9.6 222.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 222.03 -3 222.35 -2.68 ;
    END
  END ctl[37]
  PIN ctl[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 228.03 9.6 228.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 228.03 -3 228.35 -2.68 ;
    END
  END ctl[38]
  PIN ctl[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 234.03 9.6 234.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 234.03 -3 234.35 -2.68 ;
    END
  END ctl[39]
  PIN ctl[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.03 9.6 18.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 18.03 -3 18.35 -2.68 ;
    END
  END ctl[3]
  PIN ctl[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 240.03 9.6 240.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 240.03 -3 240.35 -2.68 ;
    END
  END ctl[40]
  PIN ctl[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 246.03 9.6 246.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 246.03 -3 246.35 -2.68 ;
    END
  END ctl[41]
  PIN ctl[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 252.03 9.6 252.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 252.03 -3 252.35 -2.68 ;
    END
  END ctl[42]
  PIN ctl[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 258.03 9.6 258.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 258.03 -3 258.35 -2.68 ;
    END
  END ctl[43]
  PIN ctl[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 264.03 9.6 264.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 264.03 -3 264.35 -2.68 ;
    END
  END ctl[44]
  PIN ctl[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 270.03 9.6 270.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 270.03 -3 270.35 -2.68 ;
    END
  END ctl[45]
  PIN ctl[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 276.03 9.6 276.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 276.03 -3 276.35 -2.68 ;
    END
  END ctl[46]
  PIN ctl[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 282.03 9.6 282.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 282.03 -3 282.35 -2.68 ;
    END
  END ctl[47]
  PIN ctl[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 288.03 9.6 288.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 288.03 -3 288.35 -2.68 ;
    END
  END ctl[48]
  PIN ctl[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 294.03 9.6 294.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 294.03 -3 294.35 -2.68 ;
    END
  END ctl[49]
  PIN ctl[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 24.03 9.6 24.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 24.03 -3 24.35 -2.68 ;
    END
  END ctl[4]
  PIN ctl[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 300.03 9.6 300.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 300.03 -3 300.35 -2.68 ;
    END
  END ctl[50]
  PIN ctl[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 306.03 9.6 306.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 306.03 -3 306.35 -2.68 ;
    END
  END ctl[51]
  PIN ctl[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 312.03 9.6 312.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 312.03 -3 312.35 -2.68 ;
    END
  END ctl[52]
  PIN ctl[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 318.03 9.6 318.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 318.03 -3 318.35 -2.68 ;
    END
  END ctl[53]
  PIN ctl[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 324.03 9.6 324.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 324.03 -3 324.35 -2.68 ;
    END
  END ctl[54]
  PIN ctl[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 330.03 9.6 330.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 330.03 -3 330.35 -2.68 ;
    END
  END ctl[55]
  PIN ctl[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 336.03 9.6 336.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 336.03 -3 336.35 -2.68 ;
    END
  END ctl[56]
  PIN ctl[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 342.03 9.6 342.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 342.03 -3 342.35 -2.68 ;
    END
  END ctl[57]
  PIN ctl[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 348.03 9.6 348.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 348.03 -3 348.35 -2.68 ;
    END
  END ctl[58]
  PIN ctl[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 354.03 9.6 354.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 354.03 -3 354.35 -2.68 ;
    END
  END ctl[59]
  PIN ctl[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 30.03 9.6 30.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 30.03 -3 30.35 -2.68 ;
    END
  END ctl[5]
  PIN ctl[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 360.03 9.6 360.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 360.03 -3 360.35 -2.68 ;
    END
  END ctl[60]
  PIN ctl[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 366.03 9.6 366.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 366.03 -3 366.35 -2.68 ;
    END
  END ctl[61]
  PIN ctl[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 372.03 9.6 372.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 372.03 -3 372.35 -2.68 ;
    END
  END ctl[62]
  PIN ctl[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 378.03 9.6 378.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 378.03 -3 378.35 -2.68 ;
    END
  END ctl[63]
  PIN ctl[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 384.03 9.6 384.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 384.03 -3 384.35 -2.68 ;
    END
  END ctl[64]
  PIN ctl[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 390.03 9.6 390.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 390.03 -3 390.35 -2.68 ;
    END
  END ctl[65]
  PIN ctl[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 396.03 9.6 396.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 396.03 -3 396.35 -2.68 ;
    END
  END ctl[66]
  PIN ctl[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 402.03 9.6 402.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 402.03 -3 402.35 -2.68 ;
    END
  END ctl[67]
  PIN ctl[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 408.03 9.6 408.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 408.03 -3 408.35 -2.68 ;
    END
  END ctl[68]
  PIN ctl[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 414.03 9.6 414.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 414.03 -3 414.35 -2.68 ;
    END
  END ctl[69]
  PIN ctl[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 36.03 9.6 36.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.03 -3 36.35 -2.68 ;
    END
  END ctl[6]
  PIN ctl[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 420.03 9.6 420.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 420.03 -3 420.35 -2.68 ;
    END
  END ctl[70]
  PIN ctl[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 426.03 9.6 426.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 426.03 -3 426.35 -2.68 ;
    END
  END ctl[71]
  PIN ctl[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 432.03 9.6 432.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 432.03 -3 432.35 -2.68 ;
    END
  END ctl[72]
  PIN ctl[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 438.03 9.6 438.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 438.03 -3 438.35 -2.68 ;
    END
  END ctl[73]
  PIN ctl[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 444.03 9.6 444.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 444.03 -3 444.35 -2.68 ;
    END
  END ctl[74]
  PIN ctl[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 450.03 9.6 450.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 450.03 -3 450.35 -2.68 ;
    END
  END ctl[75]
  PIN ctl[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 456.03 9.6 456.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 456.03 -3 456.35 -2.68 ;
    END
  END ctl[76]
  PIN ctl[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 462.03 9.6 462.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 462.03 -3 462.35 -2.68 ;
    END
  END ctl[77]
  PIN ctl[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 468.03 9.6 468.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 468.03 -3 468.35 -2.68 ;
    END
  END ctl[78]
  PIN ctl[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 474.03 9.6 474.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 474.03 -3 474.35 -2.68 ;
    END
  END ctl[79]
  PIN ctl[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 42.03 9.6 42.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.03 -3 42.35 -2.68 ;
    END
  END ctl[7]
  PIN ctl[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 480.03 9.6 480.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 480.03 -3 480.35 -2.68 ;
    END
  END ctl[80]
  PIN ctl[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 486.03 9.6 486.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 486.03 -3 486.35 -2.68 ;
    END
  END ctl[81]
  PIN ctl[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 492.03 9.6 492.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 492.03 -3 492.35 -2.68 ;
    END
  END ctl[82]
  PIN ctl[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 498.03 9.6 498.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 498.03 -3 498.35 -2.68 ;
    END
  END ctl[83]
  PIN ctl[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 504.03 9.6 504.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 504.03 -3 504.35 -2.68 ;
    END
  END ctl[84]
  PIN ctl[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 510.03 9.6 510.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 510.03 -3 510.35 -2.68 ;
    END
  END ctl[85]
  PIN ctl[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 516.03 9.6 516.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 516.03 -3 516.35 -2.68 ;
    END
  END ctl[86]
  PIN ctl[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 522.03 9.6 522.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 522.03 -3 522.35 -2.68 ;
    END
  END ctl[87]
  PIN ctl[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 528.03 9.6 528.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 528.03 -3 528.35 -2.68 ;
    END
  END ctl[88]
  PIN ctl[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 534.03 9.6 534.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 534.03 -3 534.35 -2.68 ;
    END
  END ctl[89]
  PIN ctl[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 48.03 9.6 48.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.03 -3 48.35 -2.68 ;
    END
  END ctl[8]
  PIN ctl[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 540.03 9.6 540.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 540.03 -3 540.35 -2.68 ;
    END
  END ctl[90]
  PIN ctl[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 546.03 9.6 546.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 546.03 -3 546.35 -2.68 ;
    END
  END ctl[91]
  PIN ctl[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 552.03 9.6 552.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 552.03 -3 552.35 -2.68 ;
    END
  END ctl[92]
  PIN ctl[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 558.03 9.6 558.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 558.03 -3 558.35 -2.68 ;
    END
  END ctl[93]
  PIN ctl[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 564.03 9.6 564.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 564.03 -3 564.35 -2.68 ;
    END
  END ctl[94]
  PIN ctl[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 570.03 9.6 570.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 570.03 -3 570.35 -2.68 ;
    END
  END ctl[95]
  PIN ctl[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 576.03 9.6 576.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 576.03 -3 576.35 -2.68 ;
    END
  END ctl[96]
  PIN ctl[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 582.03 9.6 582.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 582.03 -3 582.35 -2.68 ;
    END
  END ctl[97]
  PIN ctl[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 588.03 9.6 588.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 588.03 -3 588.35 -2.68 ;
    END
  END ctl[98]
  PIN ctl[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 594.03 9.6 594.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 594.03 -3 594.35 -2.68 ;
    END
  END ctl[99]
  PIN ctl[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 54.03 9.6 54.35 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.03 -3 54.35 -2.68 ;
    END
  END ctl[9]
  PIN ctl_b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 4.05 9.6 4.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.05 -3 4.37 -2.68 ;
    END
  END ctl_b[0]
  PIN ctl_b[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 604.05 9.6 604.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 604.05 -3 604.37 -2.68 ;
    END
  END ctl_b[100]
  PIN ctl_b[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 610.05 9.6 610.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 610.05 -3 610.37 -2.68 ;
    END
  END ctl_b[101]
  PIN ctl_b[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 616.05 9.6 616.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 616.05 -3 616.37 -2.68 ;
    END
  END ctl_b[102]
  PIN ctl_b[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 622.05 9.6 622.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 622.05 -3 622.37 -2.68 ;
    END
  END ctl_b[103]
  PIN ctl_b[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 628.05 9.6 628.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 628.05 -3 628.37 -2.68 ;
    END
  END ctl_b[104]
  PIN ctl_b[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 634.05 9.6 634.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 634.05 -3 634.37 -2.68 ;
    END
  END ctl_b[105]
  PIN ctl_b[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 640.05 9.6 640.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 640.05 -3 640.37 -2.68 ;
    END
  END ctl_b[106]
  PIN ctl_b[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 646.05 9.6 646.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 646.05 -3 646.37 -2.68 ;
    END
  END ctl_b[107]
  PIN ctl_b[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 652.05 9.6 652.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 652.05 -3 652.37 -2.68 ;
    END
  END ctl_b[108]
  PIN ctl_b[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 658.05 9.6 658.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 658.05 -3 658.37 -2.68 ;
    END
  END ctl_b[109]
  PIN ctl_b[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 64.05 9.6 64.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 64.05 -3 64.37 -2.68 ;
    END
  END ctl_b[10]
  PIN ctl_b[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 664.05 9.6 664.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 664.05 -3 664.37 -2.68 ;
    END
  END ctl_b[110]
  PIN ctl_b[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 670.05 9.6 670.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 670.05 -3 670.37 -2.68 ;
    END
  END ctl_b[111]
  PIN ctl_b[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 676.05 9.6 676.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 676.05 -3 676.37 -2.68 ;
    END
  END ctl_b[112]
  PIN ctl_b[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 682.05 9.6 682.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 682.05 -3 682.37 -2.68 ;
    END
  END ctl_b[113]
  PIN ctl_b[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 688.05 9.6 688.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 688.05 -3 688.37 -2.68 ;
    END
  END ctl_b[114]
  PIN ctl_b[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 694.05 9.6 694.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 694.05 -3 694.37 -2.68 ;
    END
  END ctl_b[115]
  PIN ctl_b[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 700.05 9.6 700.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 700.05 -3 700.37 -2.68 ;
    END
  END ctl_b[116]
  PIN ctl_b[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 706.05 9.6 706.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 706.05 -3 706.37 -2.68 ;
    END
  END ctl_b[117]
  PIN ctl_b[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 712.05 9.6 712.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 712.05 -3 712.37 -2.68 ;
    END
  END ctl_b[118]
  PIN ctl_b[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 718.05 9.6 718.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 718.05 -3 718.37 -2.68 ;
    END
  END ctl_b[119]
  PIN ctl_b[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 70.05 9.6 70.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 70.05 -3 70.37 -2.68 ;
    END
  END ctl_b[11]
  PIN ctl_b[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 724.05 9.6 724.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 724.05 -3 724.37 -2.68 ;
    END
  END ctl_b[120]
  PIN ctl_b[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 730.05 9.6 730.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 730.05 -3 730.37 -2.68 ;
    END
  END ctl_b[121]
  PIN ctl_b[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 736.05 9.6 736.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 736.05 -3 736.37 -2.68 ;
    END
  END ctl_b[122]
  PIN ctl_b[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 742.05 9.6 742.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 742.05 -3 742.37 -2.68 ;
    END
  END ctl_b[123]
  PIN ctl_b[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 748.05 9.6 748.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 748.05 -3 748.37 -2.68 ;
    END
  END ctl_b[124]
  PIN ctl_b[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 754.05 9.6 754.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 754.05 -3 754.37 -2.68 ;
    END
  END ctl_b[125]
  PIN ctl_b[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 760.05 9.6 760.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 760.05 -3 760.37 -2.68 ;
    END
  END ctl_b[126]
  PIN ctl_b[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 766.05 9.6 766.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 766.05 -3 766.37 -2.68 ;
    END
  END ctl_b[127]
  PIN ctl_b[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 76.05 9.6 76.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 76.05 -3 76.37 -2.68 ;
    END
  END ctl_b[12]
  PIN ctl_b[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 82.05 9.6 82.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.05 -3 82.37 -2.68 ;
    END
  END ctl_b[13]
  PIN ctl_b[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 88.05 9.6 88.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.05 -3 88.37 -2.68 ;
    END
  END ctl_b[14]
  PIN ctl_b[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 94.05 9.6 94.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 94.05 -3 94.37 -2.68 ;
    END
  END ctl_b[15]
  PIN ctl_b[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 100.05 9.6 100.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 100.05 -3 100.37 -2.68 ;
    END
  END ctl_b[16]
  PIN ctl_b[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 106.05 9.6 106.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 106.05 -3 106.37 -2.68 ;
    END
  END ctl_b[17]
  PIN ctl_b[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 112.05 9.6 112.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 112.05 -3 112.37 -2.68 ;
    END
  END ctl_b[18]
  PIN ctl_b[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 118.05 9.6 118.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 118.05 -3 118.37 -2.68 ;
    END
  END ctl_b[19]
  PIN ctl_b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 10.05 9.6 10.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.05 -3 10.37 -2.68 ;
    END
  END ctl_b[1]
  PIN ctl_b[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 124.05 9.6 124.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 124.05 -3 124.37 -2.68 ;
    END
  END ctl_b[20]
  PIN ctl_b[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 130.05 9.6 130.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 130.05 -3 130.37 -2.68 ;
    END
  END ctl_b[21]
  PIN ctl_b[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 136.05 9.6 136.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 136.05 -3 136.37 -2.68 ;
    END
  END ctl_b[22]
  PIN ctl_b[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 142.05 9.6 142.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 142.05 -3 142.37 -2.68 ;
    END
  END ctl_b[23]
  PIN ctl_b[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 148.05 9.6 148.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 148.05 -3 148.37 -2.68 ;
    END
  END ctl_b[24]
  PIN ctl_b[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 154.05 9.6 154.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 154.05 -3 154.37 -2.68 ;
    END
  END ctl_b[25]
  PIN ctl_b[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 160.05 9.6 160.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 160.05 -3 160.37 -2.68 ;
    END
  END ctl_b[26]
  PIN ctl_b[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 166.05 9.6 166.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 166.05 -3 166.37 -2.68 ;
    END
  END ctl_b[27]
  PIN ctl_b[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 172.05 9.6 172.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 172.05 -3 172.37 -2.68 ;
    END
  END ctl_b[28]
  PIN ctl_b[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 178.05 9.6 178.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 178.05 -3 178.37 -2.68 ;
    END
  END ctl_b[29]
  PIN ctl_b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.05 9.6 16.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 16.05 -3 16.37 -2.68 ;
    END
  END ctl_b[2]
  PIN ctl_b[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 184.05 9.6 184.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 184.05 -3 184.37 -2.68 ;
    END
  END ctl_b[30]
  PIN ctl_b[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 190.05 9.6 190.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 190.05 -3 190.37 -2.68 ;
    END
  END ctl_b[31]
  PIN ctl_b[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 196.05 9.6 196.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 196.05 -3 196.37 -2.68 ;
    END
  END ctl_b[32]
  PIN ctl_b[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 202.05 9.6 202.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 202.05 -3 202.37 -2.68 ;
    END
  END ctl_b[33]
  PIN ctl_b[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 208.05 9.6 208.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 208.05 -3 208.37 -2.68 ;
    END
  END ctl_b[34]
  PIN ctl_b[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 214.05 9.6 214.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 214.05 -3 214.37 -2.68 ;
    END
  END ctl_b[35]
  PIN ctl_b[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 220.05 9.6 220.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 220.05 -3 220.37 -2.68 ;
    END
  END ctl_b[36]
  PIN ctl_b[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 226.05 9.6 226.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 226.05 -3 226.37 -2.68 ;
    END
  END ctl_b[37]
  PIN ctl_b[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 232.05 9.6 232.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 232.05 -3 232.37 -2.68 ;
    END
  END ctl_b[38]
  PIN ctl_b[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 238.05 9.6 238.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 238.05 -3 238.37 -2.68 ;
    END
  END ctl_b[39]
  PIN ctl_b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 22.05 9.6 22.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 22.05 -3 22.37 -2.68 ;
    END
  END ctl_b[3]
  PIN ctl_b[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 244.05 9.6 244.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 244.05 -3 244.37 -2.68 ;
    END
  END ctl_b[40]
  PIN ctl_b[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 250.05 9.6 250.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 250.05 -3 250.37 -2.68 ;
    END
  END ctl_b[41]
  PIN ctl_b[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 256.05 9.6 256.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 256.05 -3 256.37 -2.68 ;
    END
  END ctl_b[42]
  PIN ctl_b[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 262.05 9.6 262.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 262.05 -3 262.37 -2.68 ;
    END
  END ctl_b[43]
  PIN ctl_b[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 268.05 9.6 268.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 268.05 -3 268.37 -2.68 ;
    END
  END ctl_b[44]
  PIN ctl_b[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 274.05 9.6 274.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 274.05 -3 274.37 -2.68 ;
    END
  END ctl_b[45]
  PIN ctl_b[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 280.05 9.6 280.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 280.05 -3 280.37 -2.68 ;
    END
  END ctl_b[46]
  PIN ctl_b[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 286.05 9.6 286.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 286.05 -3 286.37 -2.68 ;
    END
  END ctl_b[47]
  PIN ctl_b[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 292.05 9.6 292.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 292.05 -3 292.37 -2.68 ;
    END
  END ctl_b[48]
  PIN ctl_b[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 298.05 9.6 298.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 298.05 -3 298.37 -2.68 ;
    END
  END ctl_b[49]
  PIN ctl_b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 28.05 9.6 28.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 28.05 -3 28.37 -2.68 ;
    END
  END ctl_b[4]
  PIN ctl_b[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 304.05 9.6 304.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 304.05 -3 304.37 -2.68 ;
    END
  END ctl_b[50]
  PIN ctl_b[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 310.05 9.6 310.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 310.05 -3 310.37 -2.68 ;
    END
  END ctl_b[51]
  PIN ctl_b[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 316.05 9.6 316.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 316.05 -3 316.37 -2.68 ;
    END
  END ctl_b[52]
  PIN ctl_b[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 322.05 9.6 322.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 322.05 -3 322.37 -2.68 ;
    END
  END ctl_b[53]
  PIN ctl_b[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 328.05 9.6 328.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 328.05 -3 328.37 -2.68 ;
    END
  END ctl_b[54]
  PIN ctl_b[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 334.05 9.6 334.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 334.05 -3 334.37 -2.68 ;
    END
  END ctl_b[55]
  PIN ctl_b[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 340.05 9.6 340.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 340.05 -3 340.37 -2.68 ;
    END
  END ctl_b[56]
  PIN ctl_b[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 346.05 9.6 346.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 346.05 -3 346.37 -2.68 ;
    END
  END ctl_b[57]
  PIN ctl_b[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 352.05 9.6 352.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 352.05 -3 352.37 -2.68 ;
    END
  END ctl_b[58]
  PIN ctl_b[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 358.05 9.6 358.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 358.05 -3 358.37 -2.68 ;
    END
  END ctl_b[59]
  PIN ctl_b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 34.05 9.6 34.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 34.05 -3 34.37 -2.68 ;
    END
  END ctl_b[5]
  PIN ctl_b[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 364.05 9.6 364.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 364.05 -3 364.37 -2.68 ;
    END
  END ctl_b[60]
  PIN ctl_b[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 370.05 9.6 370.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 370.05 -3 370.37 -2.68 ;
    END
  END ctl_b[61]
  PIN ctl_b[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 376.05 9.6 376.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 376.05 -3 376.37 -2.68 ;
    END
  END ctl_b[62]
  PIN ctl_b[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 382.05 9.6 382.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 382.05 -3 382.37 -2.68 ;
    END
  END ctl_b[63]
  PIN ctl_b[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 388.05 9.6 388.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 388.05 -3 388.37 -2.68 ;
    END
  END ctl_b[64]
  PIN ctl_b[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 394.05 9.6 394.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 394.05 -3 394.37 -2.68 ;
    END
  END ctl_b[65]
  PIN ctl_b[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 400.05 9.6 400.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 400.05 -3 400.37 -2.68 ;
    END
  END ctl_b[66]
  PIN ctl_b[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 406.05 9.6 406.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 406.05 -3 406.37 -2.68 ;
    END
  END ctl_b[67]
  PIN ctl_b[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 412.05 9.6 412.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 412.05 -3 412.37 -2.68 ;
    END
  END ctl_b[68]
  PIN ctl_b[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 418.05 9.6 418.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 418.05 -3 418.37 -2.68 ;
    END
  END ctl_b[69]
  PIN ctl_b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 40.05 9.6 40.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 40.05 -3 40.37 -2.68 ;
    END
  END ctl_b[6]
  PIN ctl_b[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 424.05 9.6 424.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 424.05 -3 424.37 -2.68 ;
    END
  END ctl_b[70]
  PIN ctl_b[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 430.05 9.6 430.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 430.05 -3 430.37 -2.68 ;
    END
  END ctl_b[71]
  PIN ctl_b[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 436.05 9.6 436.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 436.05 -3 436.37 -2.68 ;
    END
  END ctl_b[72]
  PIN ctl_b[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 442.05 9.6 442.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 442.05 -3 442.37 -2.68 ;
    END
  END ctl_b[73]
  PIN ctl_b[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 448.05 9.6 448.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 448.05 -3 448.37 -2.68 ;
    END
  END ctl_b[74]
  PIN ctl_b[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 454.05 9.6 454.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 454.05 -3 454.37 -2.68 ;
    END
  END ctl_b[75]
  PIN ctl_b[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 460.05 9.6 460.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 460.05 -3 460.37 -2.68 ;
    END
  END ctl_b[76]
  PIN ctl_b[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 466.05 9.6 466.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 466.05 -3 466.37 -2.68 ;
    END
  END ctl_b[77]
  PIN ctl_b[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 472.05 9.6 472.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 472.05 -3 472.37 -2.68 ;
    END
  END ctl_b[78]
  PIN ctl_b[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 478.05 9.6 478.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 478.05 -3 478.37 -2.68 ;
    END
  END ctl_b[79]
  PIN ctl_b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 46.05 9.6 46.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 46.05 -3 46.37 -2.68 ;
    END
  END ctl_b[7]
  PIN ctl_b[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 484.05 9.6 484.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 484.05 -3 484.37 -2.68 ;
    END
  END ctl_b[80]
  PIN ctl_b[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 490.05 9.6 490.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 490.05 -3 490.37 -2.68 ;
    END
  END ctl_b[81]
  PIN ctl_b[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 496.05 9.6 496.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 496.05 -3 496.37 -2.68 ;
    END
  END ctl_b[82]
  PIN ctl_b[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 502.05 9.6 502.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 502.05 -3 502.37 -2.68 ;
    END
  END ctl_b[83]
  PIN ctl_b[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 508.05 9.6 508.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 508.05 -3 508.37 -2.68 ;
    END
  END ctl_b[84]
  PIN ctl_b[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 514.05 9.6 514.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 514.05 -3 514.37 -2.68 ;
    END
  END ctl_b[85]
  PIN ctl_b[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 520.05 9.6 520.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 520.05 -3 520.37 -2.68 ;
    END
  END ctl_b[86]
  PIN ctl_b[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 526.05 9.6 526.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 526.05 -3 526.37 -2.68 ;
    END
  END ctl_b[87]
  PIN ctl_b[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 532.05 9.6 532.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 532.05 -3 532.37 -2.68 ;
    END
  END ctl_b[88]
  PIN ctl_b[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 538.05 9.6 538.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 538.05 -3 538.37 -2.68 ;
    END
  END ctl_b[89]
  PIN ctl_b[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 52.05 9.6 52.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 52.05 -3 52.37 -2.68 ;
    END
  END ctl_b[8]
  PIN ctl_b[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 544.05 9.6 544.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 544.05 -3 544.37 -2.68 ;
    END
  END ctl_b[90]
  PIN ctl_b[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 550.05 9.6 550.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 550.05 -3 550.37 -2.68 ;
    END
  END ctl_b[91]
  PIN ctl_b[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 556.05 9.6 556.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 556.05 -3 556.37 -2.68 ;
    END
  END ctl_b[92]
  PIN ctl_b[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 562.05 9.6 562.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 562.05 -3 562.37 -2.68 ;
    END
  END ctl_b[93]
  PIN ctl_b[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 568.05 9.6 568.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 568.05 -3 568.37 -2.68 ;
    END
  END ctl_b[94]
  PIN ctl_b[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 574.05 9.6 574.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 574.05 -3 574.37 -2.68 ;
    END
  END ctl_b[95]
  PIN ctl_b[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 580.05 9.6 580.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 580.05 -3 580.37 -2.68 ;
    END
  END ctl_b[96]
  PIN ctl_b[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 586.05 9.6 586.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 586.05 -3 586.37 -2.68 ;
    END
  END ctl_b[97]
  PIN ctl_b[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 592.05 9.6 592.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 592.05 -3 592.37 -2.68 ;
    END
  END ctl_b[98]
  PIN ctl_b[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 598.05 9.6 598.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 598.05 -3 598.37 -2.68 ;
    END
  END ctl_b[99]
  PIN ctl_b[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 58.05 9.6 58.37 9.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 58.05 -3 58.37 -2.68 ;
    END
  END ctl_b[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 365.675 5.955 366.005 6.285 ;
        RECT 365.675 1.875 366.005 2.205 ;
        RECT 365.675 0.515 366.005 0.845 ;
        RECT 365.68 -0.16 366 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 367.035 5.955 367.365 6.285 ;
        RECT 367.035 1.875 367.365 2.205 ;
        RECT 367.035 0.515 367.365 0.845 ;
        RECT 367.04 -0.16 367.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 368.395 5.955 368.725 6.285 ;
        RECT 368.395 0.515 368.725 0.845 ;
        RECT 368.4 -0.16 368.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 369.755 5.955 370.085 6.285 ;
        RECT 369.755 0.515 370.085 0.845 ;
        RECT 369.76 -0.16 370.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 371.115 5.955 371.445 6.285 ;
        RECT 371.115 0.515 371.445 0.845 ;
        RECT 371.12 -0.16 371.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 372.475 5.955 372.805 6.285 ;
        RECT 372.475 0.515 372.805 0.845 ;
        RECT 372.48 -0.16 372.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 373.835 5.955 374.165 6.285 ;
        RECT 373.835 0.515 374.165 0.845 ;
        RECT 373.84 -0.16 374.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 375.195 5.955 375.525 6.285 ;
        RECT 375.195 0.515 375.525 0.845 ;
        RECT 375.2 -0.16 375.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 376.555 5.955 376.885 6.285 ;
        RECT 376.555 1.875 376.885 2.205 ;
        RECT 376.555 0.515 376.885 0.845 ;
        RECT 376.56 -0.16 376.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 377.915 5.955 378.245 6.285 ;
        RECT 377.915 1.875 378.245 2.205 ;
        RECT 377.915 0.515 378.245 0.845 ;
        RECT 377.92 -0.16 378.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 379.275 5.955 379.605 6.285 ;
        RECT 379.275 1.875 379.605 2.205 ;
        RECT 379.275 0.515 379.605 0.845 ;
        RECT 379.28 -0.16 379.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 380.635 5.955 380.965 6.285 ;
        RECT 380.635 0.515 380.965 0.845 ;
        RECT 380.64 -0.16 380.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 381.995 5.955 382.325 6.285 ;
        RECT 381.995 0.515 382.325 0.845 ;
        RECT 382 -0.16 382.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 383.355 5.955 383.685 6.285 ;
        RECT 383.355 0.515 383.685 0.845 ;
        RECT 383.36 -0.16 383.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 384.715 5.955 385.045 6.285 ;
        RECT 384.715 0.515 385.045 0.845 ;
        RECT 384.72 -0.16 385.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 386.075 5.955 386.405 6.285 ;
        RECT 386.075 0.515 386.405 0.845 ;
        RECT 386.08 -0.16 386.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 387.435 5.955 387.765 6.285 ;
        RECT 387.435 0.515 387.765 0.845 ;
        RECT 387.44 -0.16 387.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 388.795 5.955 389.125 6.285 ;
        RECT 388.795 1.875 389.125 2.205 ;
        RECT 388.795 0.515 389.125 0.845 ;
        RECT 388.8 -0.16 389.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 390.155 5.955 390.485 6.285 ;
        RECT 390.155 1.875 390.485 2.205 ;
        RECT 390.155 0.515 390.485 0.845 ;
        RECT 390.16 -0.16 390.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 391.515 5.955 391.845 6.285 ;
        RECT 391.515 1.875 391.845 2.205 ;
        RECT 391.515 0.515 391.845 0.845 ;
        RECT 391.52 -0.16 391.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 392.875 5.955 393.205 6.285 ;
        RECT 392.875 0.515 393.205 0.845 ;
        RECT 392.88 -0.16 393.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 394.235 5.955 394.565 6.285 ;
        RECT 394.235 0.515 394.565 0.845 ;
        RECT 394.24 -0.16 394.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 395.595 5.955 395.925 6.285 ;
        RECT 395.595 0.515 395.925 0.845 ;
        RECT 395.6 -0.16 395.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 396.955 5.955 397.285 6.285 ;
        RECT 396.955 0.515 397.285 0.845 ;
        RECT 396.96 -0.16 397.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 398.315 5.955 398.645 6.285 ;
        RECT 398.315 0.515 398.645 0.845 ;
        RECT 398.32 -0.16 398.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 399.675 5.955 400.005 6.285 ;
        RECT 399.675 1.875 400.005 2.205 ;
        RECT 399.675 0.515 400.005 0.845 ;
        RECT 399.68 -0.16 400 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 401.035 5.955 401.365 6.285 ;
        RECT 401.035 1.875 401.365 2.205 ;
        RECT 401.035 0.515 401.365 0.845 ;
        RECT 401.04 -0.16 401.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 402.395 5.955 402.725 6.285 ;
        RECT 402.395 1.875 402.725 2.205 ;
        RECT 402.395 0.515 402.725 0.845 ;
        RECT 402.4 -0.16 402.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 403.755 5.955 404.085 6.285 ;
        RECT 403.755 0.515 404.085 0.845 ;
        RECT 403.76 -0.16 404.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 405.115 5.955 405.445 6.285 ;
        RECT 405.115 0.515 405.445 0.845 ;
        RECT 405.12 -0.16 405.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 406.475 5.955 406.805 6.285 ;
        RECT 406.475 0.515 406.805 0.845 ;
        RECT 406.48 -0.16 406.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 407.835 5.955 408.165 6.285 ;
        RECT 407.835 0.515 408.165 0.845 ;
        RECT 407.84 -0.16 408.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 409.195 5.955 409.525 6.285 ;
        RECT 409.195 0.515 409.525 0.845 ;
        RECT 409.2 -0.16 409.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 410.555 5.955 410.885 6.285 ;
        RECT 410.555 0.515 410.885 0.845 ;
        RECT 410.56 -0.16 410.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 411.915 5.955 412.245 6.285 ;
        RECT 411.915 1.875 412.245 2.205 ;
        RECT 411.915 0.515 412.245 0.845 ;
        RECT 411.92 -0.16 412.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 413.275 5.955 413.605 6.285 ;
        RECT 413.275 1.875 413.605 2.205 ;
        RECT 413.275 0.515 413.605 0.845 ;
        RECT 413.28 -0.16 413.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 414.635 5.955 414.965 6.285 ;
        RECT 414.635 1.875 414.965 2.205 ;
        RECT 414.635 0.515 414.965 0.845 ;
        RECT 414.64 -0.16 414.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 415.995 5.955 416.325 6.285 ;
        RECT 415.995 0.515 416.325 0.845 ;
        RECT 416 -0.16 416.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 417.355 5.955 417.685 6.285 ;
        RECT 417.355 0.515 417.685 0.845 ;
        RECT 417.36 -0.16 417.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 418.715 5.955 419.045 6.285 ;
        RECT 418.715 0.515 419.045 0.845 ;
        RECT 418.72 -0.16 419.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 420.075 5.955 420.405 6.285 ;
        RECT 420.075 0.515 420.405 0.845 ;
        RECT 420.08 -0.16 420.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 421.435 5.955 421.765 6.285 ;
        RECT 421.435 0.515 421.765 0.845 ;
        RECT 421.44 -0.16 421.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 422.795 5.955 423.125 6.285 ;
        RECT 422.795 0.515 423.125 0.845 ;
        RECT 422.8 -0.16 423.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 424.155 5.955 424.485 6.285 ;
        RECT 424.155 1.875 424.485 2.205 ;
        RECT 424.155 0.515 424.485 0.845 ;
        RECT 424.16 -0.16 424.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 425.515 5.955 425.845 6.285 ;
        RECT 425.515 1.875 425.845 2.205 ;
        RECT 425.515 0.515 425.845 0.845 ;
        RECT 425.52 -0.16 425.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 426.875 5.955 427.205 6.285 ;
        RECT 426.875 1.875 427.205 2.205 ;
        RECT 426.875 0.515 427.205 0.845 ;
        RECT 426.88 -0.16 427.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 428.235 5.955 428.565 6.285 ;
        RECT 428.235 0.515 428.565 0.845 ;
        RECT 428.24 -0.16 428.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 429.595 5.955 429.925 6.285 ;
        RECT 429.595 0.515 429.925 0.845 ;
        RECT 429.6 -0.16 429.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 430.955 5.955 431.285 6.285 ;
        RECT 430.955 0.515 431.285 0.845 ;
        RECT 430.96 -0.16 431.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 432.315 5.955 432.645 6.285 ;
        RECT 432.315 0.515 432.645 0.845 ;
        RECT 432.32 -0.16 432.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 433.675 5.955 434.005 6.285 ;
        RECT 433.675 0.515 434.005 0.845 ;
        RECT 433.68 -0.16 434 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 435.035 5.955 435.365 6.285 ;
        RECT 435.035 0.515 435.365 0.845 ;
        RECT 435.04 -0.16 435.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 436.395 5.955 436.725 6.285 ;
        RECT 436.395 1.875 436.725 2.205 ;
        RECT 436.395 0.515 436.725 0.845 ;
        RECT 436.4 -0.16 436.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 437.755 5.955 438.085 6.285 ;
        RECT 437.755 1.875 438.085 2.205 ;
        RECT 437.755 0.515 438.085 0.845 ;
        RECT 437.76 -0.16 438.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 439.115 5.955 439.445 6.285 ;
        RECT 439.115 1.875 439.445 2.205 ;
        RECT 439.115 0.515 439.445 0.845 ;
        RECT 439.12 -0.16 439.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 440.475 5.955 440.805 6.285 ;
        RECT 440.475 0.515 440.805 0.845 ;
        RECT 440.48 -0.16 440.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 441.835 5.955 442.165 6.285 ;
        RECT 441.835 0.515 442.165 0.845 ;
        RECT 441.84 -0.16 442.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 443.195 5.955 443.525 6.285 ;
        RECT 443.195 0.515 443.525 0.845 ;
        RECT 443.2 -0.16 443.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 444.555 5.955 444.885 6.285 ;
        RECT 444.555 0.515 444.885 0.845 ;
        RECT 444.56 -0.16 444.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 445.915 5.955 446.245 6.285 ;
        RECT 445.915 0.515 446.245 0.845 ;
        RECT 445.92 -0.16 446.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 447.275 5.955 447.605 6.285 ;
        RECT 447.275 0.515 447.605 0.845 ;
        RECT 447.28 -0.16 447.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 448.635 5.955 448.965 6.285 ;
        RECT 448.635 1.875 448.965 2.205 ;
        RECT 448.635 0.515 448.965 0.845 ;
        RECT 448.64 -0.16 448.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 449.995 5.955 450.325 6.285 ;
        RECT 449.995 1.875 450.325 2.205 ;
        RECT 449.995 0.515 450.325 0.845 ;
        RECT 450 -0.16 450.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 451.355 5.955 451.685 6.285 ;
        RECT 451.355 1.875 451.685 2.205 ;
        RECT 451.355 0.515 451.685 0.845 ;
        RECT 451.36 -0.16 451.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 452.715 5.955 453.045 6.285 ;
        RECT 452.715 0.515 453.045 0.845 ;
        RECT 452.72 -0.16 453.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 454.075 5.955 454.405 6.285 ;
        RECT 454.075 0.515 454.405 0.845 ;
        RECT 454.08 -0.16 454.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 455.435 5.955 455.765 6.285 ;
        RECT 455.435 0.515 455.765 0.845 ;
        RECT 455.44 -0.16 455.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 456.795 5.955 457.125 6.285 ;
        RECT 456.795 0.515 457.125 0.845 ;
        RECT 456.8 -0.16 457.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 458.155 5.955 458.485 6.285 ;
        RECT 458.155 0.515 458.485 0.845 ;
        RECT 458.16 -0.16 458.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 459.515 5.955 459.845 6.285 ;
        RECT 459.515 1.875 459.845 2.205 ;
        RECT 459.515 0.515 459.845 0.845 ;
        RECT 459.52 -0.16 459.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 460.875 5.955 461.205 6.285 ;
        RECT 460.875 1.875 461.205 2.205 ;
        RECT 460.875 0.515 461.205 0.845 ;
        RECT 460.88 -0.16 461.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 462.235 5.955 462.565 6.285 ;
        RECT 462.235 1.875 462.565 2.205 ;
        RECT 462.235 0.515 462.565 0.845 ;
        RECT 462.24 -0.16 462.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 463.595 5.955 463.925 6.285 ;
        RECT 463.595 0.515 463.925 0.845 ;
        RECT 463.6 -0.16 463.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 464.955 5.955 465.285 6.285 ;
        RECT 464.955 0.515 465.285 0.845 ;
        RECT 464.96 -0.16 465.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 466.315 5.955 466.645 6.285 ;
        RECT 466.315 0.515 466.645 0.845 ;
        RECT 466.32 -0.16 466.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 467.675 5.955 468.005 6.285 ;
        RECT 467.675 0.515 468.005 0.845 ;
        RECT 467.68 -0.16 468 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 469.035 5.955 469.365 6.285 ;
        RECT 469.035 0.515 469.365 0.845 ;
        RECT 469.04 -0.16 469.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 470.395 5.955 470.725 6.285 ;
        RECT 470.395 0.515 470.725 0.845 ;
        RECT 470.4 -0.16 470.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 471.755 5.955 472.085 6.285 ;
        RECT 471.755 1.875 472.085 2.205 ;
        RECT 471.755 0.515 472.085 0.845 ;
        RECT 471.76 -0.16 472.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 473.115 5.955 473.445 6.285 ;
        RECT 473.115 1.875 473.445 2.205 ;
        RECT 473.115 0.515 473.445 0.845 ;
        RECT 473.12 -0.16 473.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 474.475 5.955 474.805 6.285 ;
        RECT 474.475 1.875 474.805 2.205 ;
        RECT 474.475 0.515 474.805 0.845 ;
        RECT 474.48 -0.16 474.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 475.835 5.955 476.165 6.285 ;
        RECT 475.835 0.515 476.165 0.845 ;
        RECT 475.84 -0.16 476.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 477.195 5.955 477.525 6.285 ;
        RECT 477.195 0.515 477.525 0.845 ;
        RECT 477.2 -0.16 477.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 478.555 5.955 478.885 6.285 ;
        RECT 478.555 0.515 478.885 0.845 ;
        RECT 478.56 -0.16 478.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 479.915 5.955 480.245 6.285 ;
        RECT 479.915 0.515 480.245 0.845 ;
        RECT 479.92 -0.16 480.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 481.275 5.955 481.605 6.285 ;
        RECT 481.275 0.515 481.605 0.845 ;
        RECT 481.28 -0.16 481.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 482.635 5.955 482.965 6.285 ;
        RECT 482.635 0.515 482.965 0.845 ;
        RECT 482.64 -0.16 482.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 483.995 5.955 484.325 6.285 ;
        RECT 483.995 1.875 484.325 2.205 ;
        RECT 483.995 0.515 484.325 0.845 ;
        RECT 484 -0.16 484.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 485.355 5.955 485.685 6.285 ;
        RECT 485.355 1.875 485.685 2.205 ;
        RECT 485.355 0.515 485.685 0.845 ;
        RECT 485.36 -0.16 485.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 486.715 5.955 487.045 6.285 ;
        RECT 486.715 1.875 487.045 2.205 ;
        RECT 486.715 0.515 487.045 0.845 ;
        RECT 486.72 -0.16 487.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 488.075 5.955 488.405 6.285 ;
        RECT 488.075 0.515 488.405 0.845 ;
        RECT 488.08 -0.16 488.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 489.435 5.955 489.765 6.285 ;
        RECT 489.435 0.515 489.765 0.845 ;
        RECT 489.44 -0.16 489.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 490.795 5.955 491.125 6.285 ;
        RECT 490.795 0.515 491.125 0.845 ;
        RECT 490.8 -0.16 491.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 492.155 5.955 492.485 6.285 ;
        RECT 492.155 0.515 492.485 0.845 ;
        RECT 492.16 -0.16 492.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 493.515 5.955 493.845 6.285 ;
        RECT 493.515 0.515 493.845 0.845 ;
        RECT 493.52 -0.16 493.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 494.875 5.955 495.205 6.285 ;
        RECT 494.875 0.515 495.205 0.845 ;
        RECT 494.88 -0.16 495.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 496.235 5.955 496.565 6.285 ;
        RECT 496.235 1.875 496.565 2.205 ;
        RECT 496.235 0.515 496.565 0.845 ;
        RECT 496.24 -0.16 496.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 497.595 5.955 497.925 6.285 ;
        RECT 497.595 1.875 497.925 2.205 ;
        RECT 497.595 0.515 497.925 0.845 ;
        RECT 497.6 -0.16 497.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 498.955 5.955 499.285 6.285 ;
        RECT 498.955 1.875 499.285 2.205 ;
        RECT 498.955 0.515 499.285 0.845 ;
        RECT 498.96 -0.16 499.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 500.315 5.955 500.645 6.285 ;
        RECT 500.315 0.515 500.645 0.845 ;
        RECT 500.32 -0.16 500.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 501.675 5.955 502.005 6.285 ;
        RECT 501.675 0.515 502.005 0.845 ;
        RECT 501.68 -0.16 502 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 503.035 5.955 503.365 6.285 ;
        RECT 503.035 0.515 503.365 0.845 ;
        RECT 503.04 -0.16 503.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 504.395 5.955 504.725 6.285 ;
        RECT 504.395 0.515 504.725 0.845 ;
        RECT 504.4 -0.16 504.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 505.755 5.955 506.085 6.285 ;
        RECT 505.755 0.515 506.085 0.845 ;
        RECT 505.76 -0.16 506.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 507.115 5.955 507.445 6.285 ;
        RECT 507.115 0.515 507.445 0.845 ;
        RECT 507.12 -0.16 507.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 508.475 5.955 508.805 6.285 ;
        RECT 508.475 1.875 508.805 2.205 ;
        RECT 508.475 0.515 508.805 0.845 ;
        RECT 508.48 -0.16 508.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 509.835 5.955 510.165 6.285 ;
        RECT 509.835 1.875 510.165 2.205 ;
        RECT 509.835 0.515 510.165 0.845 ;
        RECT 509.84 -0.16 510.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 511.195 5.955 511.525 6.285 ;
        RECT 511.195 1.875 511.525 2.205 ;
        RECT 511.195 0.515 511.525 0.845 ;
        RECT 511.2 -0.16 511.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 512.555 5.955 512.885 6.285 ;
        RECT 512.555 0.515 512.885 0.845 ;
        RECT 512.56 -0.16 512.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 513.915 5.955 514.245 6.285 ;
        RECT 513.915 0.515 514.245 0.845 ;
        RECT 513.92 -0.16 514.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 515.275 5.955 515.605 6.285 ;
        RECT 515.275 0.515 515.605 0.845 ;
        RECT 515.28 -0.16 515.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 516.635 5.955 516.965 6.285 ;
        RECT 516.635 0.515 516.965 0.845 ;
        RECT 516.64 -0.16 516.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 517.995 5.955 518.325 6.285 ;
        RECT 517.995 0.515 518.325 0.845 ;
        RECT 518 -0.16 518.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 519.355 5.955 519.685 6.285 ;
        RECT 519.355 0.515 519.685 0.845 ;
        RECT 519.36 -0.16 519.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 520.715 5.955 521.045 6.285 ;
        RECT 520.715 1.875 521.045 2.205 ;
        RECT 520.715 0.515 521.045 0.845 ;
        RECT 520.72 -0.16 521.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 522.075 5.955 522.405 6.285 ;
        RECT 522.075 1.875 522.405 2.205 ;
        RECT 522.075 0.515 522.405 0.845 ;
        RECT 522.08 -0.16 522.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 523.435 5.955 523.765 6.285 ;
        RECT 523.435 1.875 523.765 2.205 ;
        RECT 523.435 0.515 523.765 0.845 ;
        RECT 523.44 -0.16 523.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 524.795 5.955 525.125 6.285 ;
        RECT 524.795 0.515 525.125 0.845 ;
        RECT 524.8 -0.16 525.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 526.155 5.955 526.485 6.285 ;
        RECT 526.155 0.515 526.485 0.845 ;
        RECT 526.16 -0.16 526.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 527.515 5.955 527.845 6.285 ;
        RECT 527.515 0.515 527.845 0.845 ;
        RECT 527.52 -0.16 527.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 528.875 5.955 529.205 6.285 ;
        RECT 528.875 0.515 529.205 0.845 ;
        RECT 528.88 -0.16 529.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 530.235 5.955 530.565 6.285 ;
        RECT 530.235 0.515 530.565 0.845 ;
        RECT 530.24 -0.16 530.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 531.595 5.955 531.925 6.285 ;
        RECT 531.595 1.875 531.925 2.205 ;
        RECT 531.595 0.515 531.925 0.845 ;
        RECT 531.6 -0.16 531.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 532.955 5.955 533.285 6.285 ;
        RECT 532.955 1.875 533.285 2.205 ;
        RECT 532.955 0.515 533.285 0.845 ;
        RECT 532.96 -0.16 533.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 534.315 5.955 534.645 6.285 ;
        RECT 534.315 1.875 534.645 2.205 ;
        RECT 534.315 0.515 534.645 0.845 ;
        RECT 534.32 -0.16 534.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 535.675 5.955 536.005 6.285 ;
        RECT 535.675 0.515 536.005 0.845 ;
        RECT 535.68 -0.16 536 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 537.035 5.955 537.365 6.285 ;
        RECT 537.035 0.515 537.365 0.845 ;
        RECT 537.04 -0.16 537.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 538.395 5.955 538.725 6.285 ;
        RECT 538.395 0.515 538.725 0.845 ;
        RECT 538.4 -0.16 538.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 539.755 5.955 540.085 6.285 ;
        RECT 539.755 0.515 540.085 0.845 ;
        RECT 539.76 -0.16 540.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 541.115 5.955 541.445 6.285 ;
        RECT 541.115 0.515 541.445 0.845 ;
        RECT 541.12 -0.16 541.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 542.475 5.955 542.805 6.285 ;
        RECT 542.475 0.515 542.805 0.845 ;
        RECT 542.48 -0.16 542.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 543.835 5.955 544.165 6.285 ;
        RECT 543.835 1.875 544.165 2.205 ;
        RECT 543.835 0.515 544.165 0.845 ;
        RECT 543.84 -0.16 544.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 545.195 5.955 545.525 6.285 ;
        RECT 545.195 1.875 545.525 2.205 ;
        RECT 545.195 0.515 545.525 0.845 ;
        RECT 545.2 -0.16 545.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 546.555 5.955 546.885 6.285 ;
        RECT 546.555 1.875 546.885 2.205 ;
        RECT 546.555 0.515 546.885 0.845 ;
        RECT 546.56 -0.16 546.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 547.915 5.955 548.245 6.285 ;
        RECT 547.915 0.515 548.245 0.845 ;
        RECT 547.92 -0.16 548.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 549.275 5.955 549.605 6.285 ;
        RECT 549.275 0.515 549.605 0.845 ;
        RECT 549.28 -0.16 549.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 550.635 5.955 550.965 6.285 ;
        RECT 550.635 0.515 550.965 0.845 ;
        RECT 550.64 -0.16 550.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 551.995 5.955 552.325 6.285 ;
        RECT 551.995 0.515 552.325 0.845 ;
        RECT 552 -0.16 552.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 553.355 5.955 553.685 6.285 ;
        RECT 553.355 0.515 553.685 0.845 ;
        RECT 553.36 -0.16 553.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 554.715 5.955 555.045 6.285 ;
        RECT 554.715 0.515 555.045 0.845 ;
        RECT 554.72 -0.16 555.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 556.075 5.955 556.405 6.285 ;
        RECT 556.075 1.875 556.405 2.205 ;
        RECT 556.075 0.515 556.405 0.845 ;
        RECT 556.08 -0.16 556.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 557.435 5.955 557.765 6.285 ;
        RECT 557.435 1.875 557.765 2.205 ;
        RECT 557.435 0.515 557.765 0.845 ;
        RECT 557.44 -0.16 557.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 558.795 5.955 559.125 6.285 ;
        RECT 558.795 1.875 559.125 2.205 ;
        RECT 558.795 0.515 559.125 0.845 ;
        RECT 558.8 -0.16 559.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 560.155 5.955 560.485 6.285 ;
        RECT 560.155 0.515 560.485 0.845 ;
        RECT 560.16 -0.16 560.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 561.515 5.955 561.845 6.285 ;
        RECT 561.515 0.515 561.845 0.845 ;
        RECT 561.52 -0.16 561.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 562.875 5.955 563.205 6.285 ;
        RECT 562.875 0.515 563.205 0.845 ;
        RECT 562.88 -0.16 563.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 564.235 5.955 564.565 6.285 ;
        RECT 564.235 0.515 564.565 0.845 ;
        RECT 564.24 -0.16 564.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 565.595 5.955 565.925 6.285 ;
        RECT 565.595 0.515 565.925 0.845 ;
        RECT 565.6 -0.16 565.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 566.955 5.955 567.285 6.285 ;
        RECT 566.955 0.515 567.285 0.845 ;
        RECT 566.96 -0.16 567.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 568.315 5.955 568.645 6.285 ;
        RECT 568.315 1.875 568.645 2.205 ;
        RECT 568.315 0.515 568.645 0.845 ;
        RECT 568.32 -0.16 568.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 569.675 5.955 570.005 6.285 ;
        RECT 569.675 1.875 570.005 2.205 ;
        RECT 569.675 0.515 570.005 0.845 ;
        RECT 569.68 -0.16 570 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 571.035 5.955 571.365 6.285 ;
        RECT 571.035 1.875 571.365 2.205 ;
        RECT 571.035 0.515 571.365 0.845 ;
        RECT 571.04 -0.16 571.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 572.395 5.955 572.725 6.285 ;
        RECT 572.395 0.515 572.725 0.845 ;
        RECT 572.4 -0.16 572.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 573.755 5.955 574.085 6.285 ;
        RECT 573.755 0.515 574.085 0.845 ;
        RECT 573.76 -0.16 574.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 575.115 5.955 575.445 6.285 ;
        RECT 575.115 0.515 575.445 0.845 ;
        RECT 575.12 -0.16 575.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 576.475 5.955 576.805 6.285 ;
        RECT 576.475 0.515 576.805 0.845 ;
        RECT 576.48 -0.16 576.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 577.835 5.955 578.165 6.285 ;
        RECT 577.835 0.515 578.165 0.845 ;
        RECT 577.84 -0.16 578.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 579.195 5.955 579.525 6.285 ;
        RECT 579.195 0.515 579.525 0.845 ;
        RECT 579.2 -0.16 579.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 580.555 5.955 580.885 6.285 ;
        RECT 580.555 1.875 580.885 2.205 ;
        RECT 580.555 0.515 580.885 0.845 ;
        RECT 580.56 -0.16 580.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 581.915 5.955 582.245 6.285 ;
        RECT 581.915 1.875 582.245 2.205 ;
        RECT 581.915 0.515 582.245 0.845 ;
        RECT 581.92 -0.16 582.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 583.275 5.955 583.605 6.285 ;
        RECT 583.275 1.875 583.605 2.205 ;
        RECT 583.275 0.515 583.605 0.845 ;
        RECT 583.28 -0.16 583.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 584.635 5.955 584.965 6.285 ;
        RECT 584.635 0.515 584.965 0.845 ;
        RECT 584.64 -0.16 584.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 585.995 5.955 586.325 6.285 ;
        RECT 585.995 0.515 586.325 0.845 ;
        RECT 586 -0.16 586.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 587.355 5.955 587.685 6.285 ;
        RECT 587.355 0.515 587.685 0.845 ;
        RECT 587.36 -0.16 587.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 588.715 5.955 589.045 6.285 ;
        RECT 588.715 0.515 589.045 0.845 ;
        RECT 588.72 -0.16 589.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 590.075 5.955 590.405 6.285 ;
        RECT 590.075 0.515 590.405 0.845 ;
        RECT 590.08 -0.16 590.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 591.435 5.955 591.765 6.285 ;
        RECT 591.435 0.515 591.765 0.845 ;
        RECT 591.44 -0.16 591.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 592.795 5.955 593.125 6.285 ;
        RECT 592.795 1.875 593.125 2.205 ;
        RECT 592.795 0.515 593.125 0.845 ;
        RECT 592.8 -0.16 593.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 594.155 5.955 594.485 6.285 ;
        RECT 594.155 1.875 594.485 2.205 ;
        RECT 594.155 0.515 594.485 0.845 ;
        RECT 594.16 -0.16 594.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 595.515 5.955 595.845 6.285 ;
        RECT 595.515 1.875 595.845 2.205 ;
        RECT 595.515 0.515 595.845 0.845 ;
        RECT 595.52 -0.16 595.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 596.875 5.955 597.205 6.285 ;
        RECT 596.875 0.515 597.205 0.845 ;
        RECT 596.88 -0.16 597.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 598.235 5.955 598.565 6.285 ;
        RECT 598.235 0.515 598.565 0.845 ;
        RECT 598.24 -0.16 598.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 599.595 5.955 599.925 6.285 ;
        RECT 599.595 0.515 599.925 0.845 ;
        RECT 599.6 -0.16 599.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 600.955 5.955 601.285 6.285 ;
        RECT 600.955 0.515 601.285 0.845 ;
        RECT 600.96 -0.16 601.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 602.315 5.955 602.645 6.285 ;
        RECT 602.315 0.515 602.645 0.845 ;
        RECT 602.32 -0.16 602.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 603.675 5.955 604.005 6.285 ;
        RECT 603.675 1.875 604.005 2.205 ;
        RECT 603.675 0.515 604.005 0.845 ;
        RECT 603.68 -0.16 604 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 605.035 5.955 605.365 6.285 ;
        RECT 605.035 1.875 605.365 2.205 ;
        RECT 605.035 0.515 605.365 0.845 ;
        RECT 605.04 -0.16 605.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 606.395 5.955 606.725 6.285 ;
        RECT 606.395 1.875 606.725 2.205 ;
        RECT 606.395 0.515 606.725 0.845 ;
        RECT 606.4 -0.16 606.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 607.755 5.955 608.085 6.285 ;
        RECT 607.755 0.515 608.085 0.845 ;
        RECT 607.76 -0.16 608.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 609.115 5.955 609.445 6.285 ;
        RECT 609.115 0.515 609.445 0.845 ;
        RECT 609.12 -0.16 609.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 610.475 5.955 610.805 6.285 ;
        RECT 610.475 0.515 610.805 0.845 ;
        RECT 610.48 -0.16 610.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 611.835 5.955 612.165 6.285 ;
        RECT 611.835 0.515 612.165 0.845 ;
        RECT 611.84 -0.16 612.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 613.195 5.955 613.525 6.285 ;
        RECT 613.195 0.515 613.525 0.845 ;
        RECT 613.2 -0.16 613.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 614.555 5.955 614.885 6.285 ;
        RECT 614.555 0.515 614.885 0.845 ;
        RECT 614.56 -0.16 614.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 615.915 5.955 616.245 6.285 ;
        RECT 615.915 1.875 616.245 2.205 ;
        RECT 615.915 0.515 616.245 0.845 ;
        RECT 615.92 -0.16 616.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 617.275 5.955 617.605 6.285 ;
        RECT 617.275 1.875 617.605 2.205 ;
        RECT 617.275 0.515 617.605 0.845 ;
        RECT 617.28 -0.16 617.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 618.635 5.955 618.965 6.285 ;
        RECT 618.635 1.875 618.965 2.205 ;
        RECT 618.635 0.515 618.965 0.845 ;
        RECT 618.64 -0.16 618.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 619.995 5.955 620.325 6.285 ;
        RECT 619.995 0.515 620.325 0.845 ;
        RECT 620 -0.16 620.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 621.355 5.955 621.685 6.285 ;
        RECT 621.355 0.515 621.685 0.845 ;
        RECT 621.36 -0.16 621.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 622.715 5.955 623.045 6.285 ;
        RECT 622.715 0.515 623.045 0.845 ;
        RECT 622.72 -0.16 623.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 624.075 5.955 624.405 6.285 ;
        RECT 624.075 0.515 624.405 0.845 ;
        RECT 624.08 -0.16 624.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 625.435 5.955 625.765 6.285 ;
        RECT 625.435 0.515 625.765 0.845 ;
        RECT 625.44 -0.16 625.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 626.795 5.955 627.125 6.285 ;
        RECT 626.795 0.515 627.125 0.845 ;
        RECT 626.8 -0.16 627.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 628.155 5.955 628.485 6.285 ;
        RECT 628.155 1.875 628.485 2.205 ;
        RECT 628.155 0.515 628.485 0.845 ;
        RECT 628.16 -0.16 628.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 629.515 5.955 629.845 6.285 ;
        RECT 629.515 1.875 629.845 2.205 ;
        RECT 629.515 0.515 629.845 0.845 ;
        RECT 629.52 -0.16 629.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 630.875 5.955 631.205 6.285 ;
        RECT 630.875 1.875 631.205 2.205 ;
        RECT 630.875 0.515 631.205 0.845 ;
        RECT 630.88 -0.16 631.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 632.235 5.955 632.565 6.285 ;
        RECT 632.235 0.515 632.565 0.845 ;
        RECT 632.24 -0.16 632.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 633.595 5.955 633.925 6.285 ;
        RECT 633.595 0.515 633.925 0.845 ;
        RECT 633.6 -0.16 633.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 634.955 5.955 635.285 6.285 ;
        RECT 634.955 0.515 635.285 0.845 ;
        RECT 634.96 -0.16 635.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 636.315 5.955 636.645 6.285 ;
        RECT 636.315 0.515 636.645 0.845 ;
        RECT 636.32 -0.16 636.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 637.675 5.955 638.005 6.285 ;
        RECT 637.675 0.515 638.005 0.845 ;
        RECT 637.68 -0.16 638 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 639.035 5.955 639.365 6.285 ;
        RECT 639.035 0.515 639.365 0.845 ;
        RECT 639.04 -0.16 639.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 640.395 5.955 640.725 6.285 ;
        RECT 640.395 1.875 640.725 2.205 ;
        RECT 640.395 0.515 640.725 0.845 ;
        RECT 640.4 -0.16 640.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 641.755 5.955 642.085 6.285 ;
        RECT 641.755 1.875 642.085 2.205 ;
        RECT 641.755 0.515 642.085 0.845 ;
        RECT 641.76 -0.16 642.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 643.115 5.955 643.445 6.285 ;
        RECT 643.115 1.875 643.445 2.205 ;
        RECT 643.115 0.515 643.445 0.845 ;
        RECT 643.12 -0.16 643.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 644.475 5.955 644.805 6.285 ;
        RECT 644.475 0.515 644.805 0.845 ;
        RECT 644.48 -0.16 644.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 645.835 5.955 646.165 6.285 ;
        RECT 645.835 0.515 646.165 0.845 ;
        RECT 645.84 -0.16 646.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 647.195 5.955 647.525 6.285 ;
        RECT 647.195 0.515 647.525 0.845 ;
        RECT 647.2 -0.16 647.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 648.555 5.955 648.885 6.285 ;
        RECT 648.555 0.515 648.885 0.845 ;
        RECT 648.56 -0.16 648.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 649.915 5.955 650.245 6.285 ;
        RECT 649.915 0.515 650.245 0.845 ;
        RECT 649.92 -0.16 650.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 651.275 5.955 651.605 6.285 ;
        RECT 651.275 0.515 651.605 0.845 ;
        RECT 651.28 -0.16 651.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 652.635 5.955 652.965 6.285 ;
        RECT 652.635 1.875 652.965 2.205 ;
        RECT 652.635 0.515 652.965 0.845 ;
        RECT 652.64 -0.16 652.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 653.995 5.955 654.325 6.285 ;
        RECT 653.995 1.875 654.325 2.205 ;
        RECT 653.995 0.515 654.325 0.845 ;
        RECT 654 -0.16 654.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 655.355 5.955 655.685 6.285 ;
        RECT 655.355 1.875 655.685 2.205 ;
        RECT 655.355 0.515 655.685 0.845 ;
        RECT 655.36 -0.16 655.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 656.715 5.955 657.045 6.285 ;
        RECT 656.715 0.515 657.045 0.845 ;
        RECT 656.72 -0.16 657.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 658.075 5.955 658.405 6.285 ;
        RECT 658.075 0.515 658.405 0.845 ;
        RECT 658.08 -0.16 658.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 659.435 5.955 659.765 6.285 ;
        RECT 659.435 0.515 659.765 0.845 ;
        RECT 659.44 -0.16 659.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 660.795 5.955 661.125 6.285 ;
        RECT 660.795 0.515 661.125 0.845 ;
        RECT 660.8 -0.16 661.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 662.155 5.955 662.485 6.285 ;
        RECT 662.155 0.515 662.485 0.845 ;
        RECT 662.16 -0.16 662.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 663.515 5.955 663.845 6.285 ;
        RECT 663.515 1.875 663.845 2.205 ;
        RECT 663.515 0.515 663.845 0.845 ;
        RECT 663.52 -0.16 663.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 664.875 5.955 665.205 6.285 ;
        RECT 664.875 1.875 665.205 2.205 ;
        RECT 664.875 0.515 665.205 0.845 ;
        RECT 664.88 -0.16 665.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 666.235 5.955 666.565 6.285 ;
        RECT 666.235 1.875 666.565 2.205 ;
        RECT 666.235 0.515 666.565 0.845 ;
        RECT 666.24 -0.16 666.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 667.595 5.955 667.925 6.285 ;
        RECT 667.595 0.515 667.925 0.845 ;
        RECT 667.6 -0.16 667.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 668.955 5.955 669.285 6.285 ;
        RECT 668.955 0.515 669.285 0.845 ;
        RECT 668.96 -0.16 669.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 670.315 5.955 670.645 6.285 ;
        RECT 670.315 0.515 670.645 0.845 ;
        RECT 670.32 -0.16 670.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 671.675 5.955 672.005 6.285 ;
        RECT 671.675 0.515 672.005 0.845 ;
        RECT 671.68 -0.16 672 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 673.035 5.955 673.365 6.285 ;
        RECT 673.035 0.515 673.365 0.845 ;
        RECT 673.04 -0.16 673.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 674.395 5.955 674.725 6.285 ;
        RECT 674.395 0.515 674.725 0.845 ;
        RECT 674.4 -0.16 674.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 675.755 5.955 676.085 6.285 ;
        RECT 675.755 1.875 676.085 2.205 ;
        RECT 675.755 0.515 676.085 0.845 ;
        RECT 675.76 -0.16 676.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 677.115 5.955 677.445 6.285 ;
        RECT 677.115 1.875 677.445 2.205 ;
        RECT 677.115 0.515 677.445 0.845 ;
        RECT 677.12 -0.16 677.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 678.475 5.955 678.805 6.285 ;
        RECT 678.475 1.875 678.805 2.205 ;
        RECT 678.475 0.515 678.805 0.845 ;
        RECT 678.48 -0.16 678.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 679.835 5.955 680.165 6.285 ;
        RECT 679.835 0.515 680.165 0.845 ;
        RECT 679.84 -0.16 680.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 681.195 5.955 681.525 6.285 ;
        RECT 681.195 0.515 681.525 0.845 ;
        RECT 681.2 -0.16 681.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 682.555 5.955 682.885 6.285 ;
        RECT 682.555 0.515 682.885 0.845 ;
        RECT 682.56 -0.16 682.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 683.915 5.955 684.245 6.285 ;
        RECT 683.915 0.515 684.245 0.845 ;
        RECT 683.92 -0.16 684.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 685.275 5.955 685.605 6.285 ;
        RECT 685.275 0.515 685.605 0.845 ;
        RECT 685.28 -0.16 685.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 686.635 5.955 686.965 6.285 ;
        RECT 686.635 0.515 686.965 0.845 ;
        RECT 686.64 -0.16 686.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 687.995 5.955 688.325 6.285 ;
        RECT 687.995 1.875 688.325 2.205 ;
        RECT 687.995 0.515 688.325 0.845 ;
        RECT 688 -0.16 688.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 689.355 5.955 689.685 6.285 ;
        RECT 689.355 1.875 689.685 2.205 ;
        RECT 689.355 0.515 689.685 0.845 ;
        RECT 689.36 -0.16 689.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 690.715 5.955 691.045 6.285 ;
        RECT 690.715 1.875 691.045 2.205 ;
        RECT 690.715 0.515 691.045 0.845 ;
        RECT 690.72 -0.16 691.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 692.075 5.955 692.405 6.285 ;
        RECT 692.075 0.515 692.405 0.845 ;
        RECT 692.08 -0.16 692.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 693.435 5.955 693.765 6.285 ;
        RECT 693.435 0.515 693.765 0.845 ;
        RECT 693.44 -0.16 693.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 694.795 5.955 695.125 6.285 ;
        RECT 694.795 0.515 695.125 0.845 ;
        RECT 694.8 -0.16 695.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 696.155 5.955 696.485 6.285 ;
        RECT 696.155 0.515 696.485 0.845 ;
        RECT 696.16 -0.16 696.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 697.515 5.955 697.845 6.285 ;
        RECT 697.515 0.515 697.845 0.845 ;
        RECT 697.52 -0.16 697.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 698.875 5.955 699.205 6.285 ;
        RECT 698.875 0.515 699.205 0.845 ;
        RECT 698.88 -0.16 699.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 700.235 5.955 700.565 6.285 ;
        RECT 700.235 1.875 700.565 2.205 ;
        RECT 700.235 0.515 700.565 0.845 ;
        RECT 700.24 -0.16 700.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 701.595 5.955 701.925 6.285 ;
        RECT 701.595 1.875 701.925 2.205 ;
        RECT 701.595 0.515 701.925 0.845 ;
        RECT 701.6 -0.16 701.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 702.955 5.955 703.285 6.285 ;
        RECT 702.955 1.875 703.285 2.205 ;
        RECT 702.955 0.515 703.285 0.845 ;
        RECT 702.96 -0.16 703.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 704.315 5.955 704.645 6.285 ;
        RECT 704.315 0.515 704.645 0.845 ;
        RECT 704.32 -0.16 704.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 705.675 5.955 706.005 6.285 ;
        RECT 705.675 0.515 706.005 0.845 ;
        RECT 705.68 -0.16 706 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 707.035 5.955 707.365 6.285 ;
        RECT 707.035 0.515 707.365 0.845 ;
        RECT 707.04 -0.16 707.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 708.395 5.955 708.725 6.285 ;
        RECT 708.395 0.515 708.725 0.845 ;
        RECT 708.4 -0.16 708.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 709.755 5.955 710.085 6.285 ;
        RECT 709.755 0.515 710.085 0.845 ;
        RECT 709.76 -0.16 710.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 711.115 5.955 711.445 6.285 ;
        RECT 711.115 0.515 711.445 0.845 ;
        RECT 711.12 -0.16 711.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 712.475 5.955 712.805 6.285 ;
        RECT 712.475 1.875 712.805 2.205 ;
        RECT 712.475 0.515 712.805 0.845 ;
        RECT 712.48 -0.16 712.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 713.835 5.955 714.165 6.285 ;
        RECT 713.835 1.875 714.165 2.205 ;
        RECT 713.835 0.515 714.165 0.845 ;
        RECT 713.84 -0.16 714.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 715.195 5.955 715.525 6.285 ;
        RECT 715.195 1.875 715.525 2.205 ;
        RECT 715.195 0.515 715.525 0.845 ;
        RECT 715.2 -0.16 715.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 716.555 5.955 716.885 6.285 ;
        RECT 716.555 0.515 716.885 0.845 ;
        RECT 716.56 -0.16 716.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 717.915 5.955 718.245 6.285 ;
        RECT 717.915 0.515 718.245 0.845 ;
        RECT 717.92 -0.16 718.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 719.275 5.955 719.605 6.285 ;
        RECT 719.275 0.515 719.605 0.845 ;
        RECT 719.28 -0.16 719.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 720.635 5.955 720.965 6.285 ;
        RECT 720.635 0.515 720.965 0.845 ;
        RECT 720.64 -0.16 720.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 721.995 5.955 722.325 6.285 ;
        RECT 721.995 0.515 722.325 0.845 ;
        RECT 722 -0.16 722.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 723.355 5.955 723.685 6.285 ;
        RECT 723.355 0.515 723.685 0.845 ;
        RECT 723.36 -0.16 723.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 724.715 5.955 725.045 6.285 ;
        RECT 724.715 1.875 725.045 2.205 ;
        RECT 724.715 0.515 725.045 0.845 ;
        RECT 724.72 -0.16 725.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 726.075 5.955 726.405 6.285 ;
        RECT 726.075 1.875 726.405 2.205 ;
        RECT 726.075 0.515 726.405 0.845 ;
        RECT 726.08 -0.16 726.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 727.435 5.955 727.765 6.285 ;
        RECT 727.435 1.875 727.765 2.205 ;
        RECT 727.435 0.515 727.765 0.845 ;
        RECT 727.44 -0.16 727.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 728.795 5.955 729.125 6.285 ;
        RECT 728.795 0.515 729.125 0.845 ;
        RECT 728.8 -0.16 729.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 730.155 5.955 730.485 6.285 ;
        RECT 730.155 0.515 730.485 0.845 ;
        RECT 730.16 -0.16 730.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 731.515 5.955 731.845 6.285 ;
        RECT 731.515 0.515 731.845 0.845 ;
        RECT 731.52 -0.16 731.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 732.875 5.955 733.205 6.285 ;
        RECT 732.875 0.515 733.205 0.845 ;
        RECT 732.88 -0.16 733.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 734.235 5.955 734.565 6.285 ;
        RECT 734.235 0.515 734.565 0.845 ;
        RECT 734.24 -0.16 734.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 735.595 5.955 735.925 6.285 ;
        RECT 735.595 1.875 735.925 2.205 ;
        RECT 735.595 0.515 735.925 0.845 ;
        RECT 735.6 -0.16 735.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 736.955 5.955 737.285 6.285 ;
        RECT 736.955 1.875 737.285 2.205 ;
        RECT 736.955 0.515 737.285 0.845 ;
        RECT 736.96 -0.16 737.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 738.315 5.955 738.645 6.285 ;
        RECT 738.315 1.875 738.645 2.205 ;
        RECT 738.315 0.515 738.645 0.845 ;
        RECT 738.32 -0.16 738.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 739.675 5.955 740.005 6.285 ;
        RECT 739.675 0.515 740.005 0.845 ;
        RECT 739.68 -0.16 740 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 741.035 5.955 741.365 6.285 ;
        RECT 741.035 0.515 741.365 0.845 ;
        RECT 741.04 -0.16 741.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 742.395 5.955 742.725 6.285 ;
        RECT 742.395 0.515 742.725 0.845 ;
        RECT 742.4 -0.16 742.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 743.755 5.955 744.085 6.285 ;
        RECT 743.755 0.515 744.085 0.845 ;
        RECT 743.76 -0.16 744.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 745.115 5.955 745.445 6.285 ;
        RECT 745.115 0.515 745.445 0.845 ;
        RECT 745.12 -0.16 745.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 746.475 5.955 746.805 6.285 ;
        RECT 746.475 0.515 746.805 0.845 ;
        RECT 746.48 -0.16 746.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 747.835 5.955 748.165 6.285 ;
        RECT 747.835 1.875 748.165 2.205 ;
        RECT 747.835 0.515 748.165 0.845 ;
        RECT 747.84 -0.16 748.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 749.195 5.955 749.525 6.285 ;
        RECT 749.195 1.875 749.525 2.205 ;
        RECT 749.195 0.515 749.525 0.845 ;
        RECT 749.2 -0.16 749.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 750.555 5.955 750.885 6.285 ;
        RECT 750.555 1.875 750.885 2.205 ;
        RECT 750.555 0.515 750.885 0.845 ;
        RECT 750.56 -0.16 750.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 751.915 5.955 752.245 6.285 ;
        RECT 751.915 0.515 752.245 0.845 ;
        RECT 751.92 -0.16 752.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 753.275 5.955 753.605 6.285 ;
        RECT 753.275 0.515 753.605 0.845 ;
        RECT 753.28 -0.16 753.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 754.635 5.955 754.965 6.285 ;
        RECT 754.635 0.515 754.965 0.845 ;
        RECT 754.64 -0.16 754.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 755.995 5.955 756.325 6.285 ;
        RECT 755.995 0.515 756.325 0.845 ;
        RECT 756 -0.16 756.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 757.355 5.955 757.685 6.285 ;
        RECT 757.355 0.515 757.685 0.845 ;
        RECT 757.36 -0.16 757.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 758.715 5.955 759.045 6.285 ;
        RECT 758.715 0.515 759.045 0.845 ;
        RECT 758.72 -0.16 759.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 760.075 5.955 760.405 6.285 ;
        RECT 760.075 1.875 760.405 2.205 ;
        RECT 760.075 0.515 760.405 0.845 ;
        RECT 760.08 -0.16 760.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 761.435 5.955 761.765 6.285 ;
        RECT 761.435 1.875 761.765 2.205 ;
        RECT 761.435 0.515 761.765 0.845 ;
        RECT 761.44 -0.16 761.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 762.795 5.955 763.125 6.285 ;
        RECT 762.795 1.875 763.125 2.205 ;
        RECT 762.795 0.515 763.125 0.845 ;
        RECT 762.8 -0.16 763.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 764.155 5.955 764.485 6.285 ;
        RECT 764.155 1.875 764.485 2.205 ;
        RECT 764.155 0.515 764.485 0.845 ;
        RECT 764.16 -0.16 764.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 765.515 5.955 765.845 6.285 ;
        RECT 765.515 3.235 765.845 3.565 ;
        RECT 765.515 1.875 765.845 2.205 ;
        RECT 765.515 0.515 765.845 0.845 ;
        RECT 765.52 -0.16 765.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 766.875 5.955 767.205 6.285 ;
        RECT 766.875 3.235 767.205 3.565 ;
        RECT 766.875 1.875 767.205 2.205 ;
        RECT 766.875 0.515 767.205 0.845 ;
        RECT 766.88 -0.16 767.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 768.235 5.955 768.565 6.285 ;
        RECT 768.235 4.595 768.565 4.925 ;
        RECT 768.235 3.235 768.565 3.565 ;
        RECT 768.235 1.875 768.565 2.205 ;
        RECT 768.235 0.515 768.565 0.845 ;
        RECT 768.24 -0.16 768.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.525 5.955 -1.195 6.285 ;
        RECT -1.525 4.595 -1.195 4.925 ;
        RECT -1.525 3.235 -1.195 3.565 ;
        RECT -1.525 1.875 -1.195 2.205 ;
        RECT -1.525 0.515 -1.195 0.845 ;
        RECT -1.52 -0.16 -1.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.165 5.955 0.165 6.285 ;
        RECT -0.165 4.595 0.165 4.925 ;
        RECT -0.165 3.235 0.165 3.565 ;
        RECT -0.165 1.875 0.165 2.205 ;
        RECT -0.165 0.515 0.165 0.845 ;
        RECT -0.16 -0.16 0.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.195 5.955 1.525 6.285 ;
        RECT 1.195 3.235 1.525 3.565 ;
        RECT 1.195 1.875 1.525 2.205 ;
        RECT 1.195 0.515 1.525 0.845 ;
        RECT 1.2 -0.16 1.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 5.955 2.885 6.285 ;
        RECT 2.555 1.875 2.885 2.205 ;
        RECT 2.555 0.515 2.885 0.845 ;
        RECT 2.56 -0.16 2.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.915 5.955 4.245 6.285 ;
        RECT 3.915 1.875 4.245 2.205 ;
        RECT 3.915 0.515 4.245 0.845 ;
        RECT 3.92 -0.16 4.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.275 5.955 5.605 6.285 ;
        RECT 5.275 1.875 5.605 2.205 ;
        RECT 5.275 0.515 5.605 0.845 ;
        RECT 5.28 -0.16 5.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 5.955 6.965 6.285 ;
        RECT 6.635 1.875 6.965 2.205 ;
        RECT 6.635 0.515 6.965 0.845 ;
        RECT 6.64 -0.16 6.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.995 5.955 8.325 6.285 ;
        RECT 7.995 0.515 8.325 0.845 ;
        RECT 8 -0.16 8.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 5.955 9.685 6.285 ;
        RECT 9.355 0.515 9.685 0.845 ;
        RECT 9.36 -0.16 9.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.715 5.955 11.045 6.285 ;
        RECT 10.715 0.515 11.045 0.845 ;
        RECT 10.72 -0.16 11.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.075 5.955 12.405 6.285 ;
        RECT 12.075 0.515 12.405 0.845 ;
        RECT 12.08 -0.16 12.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.435 5.955 13.765 6.285 ;
        RECT 13.435 0.515 13.765 0.845 ;
        RECT 13.44 -0.16 13.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.795 5.955 15.125 6.285 ;
        RECT 14.795 0.515 15.125 0.845 ;
        RECT 14.8 -0.16 15.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.155 5.955 16.485 6.285 ;
        RECT 16.155 1.875 16.485 2.205 ;
        RECT 16.155 0.515 16.485 0.845 ;
        RECT 16.16 -0.16 16.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.515 5.955 17.845 6.285 ;
        RECT 17.515 1.875 17.845 2.205 ;
        RECT 17.515 0.515 17.845 0.845 ;
        RECT 17.52 -0.16 17.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.875 5.955 19.205 6.285 ;
        RECT 18.875 1.875 19.205 2.205 ;
        RECT 18.875 0.515 19.205 0.845 ;
        RECT 18.88 -0.16 19.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.235 5.955 20.565 6.285 ;
        RECT 20.235 0.515 20.565 0.845 ;
        RECT 20.24 -0.16 20.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.595 5.955 21.925 6.285 ;
        RECT 21.595 0.515 21.925 0.845 ;
        RECT 21.6 -0.16 21.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.955 5.955 23.285 6.285 ;
        RECT 22.955 0.515 23.285 0.845 ;
        RECT 22.96 -0.16 23.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.315 5.955 24.645 6.285 ;
        RECT 24.315 0.515 24.645 0.845 ;
        RECT 24.32 -0.16 24.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.675 5.955 26.005 6.285 ;
        RECT 25.675 0.515 26.005 0.845 ;
        RECT 25.68 -0.16 26 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.035 5.955 27.365 6.285 ;
        RECT 27.035 0.515 27.365 0.845 ;
        RECT 27.04 -0.16 27.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.395 5.955 28.725 6.285 ;
        RECT 28.395 1.875 28.725 2.205 ;
        RECT 28.395 0.515 28.725 0.845 ;
        RECT 28.4 -0.16 28.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.755 5.955 30.085 6.285 ;
        RECT 29.755 1.875 30.085 2.205 ;
        RECT 29.755 0.515 30.085 0.845 ;
        RECT 29.76 -0.16 30.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.115 5.955 31.445 6.285 ;
        RECT 31.115 1.875 31.445 2.205 ;
        RECT 31.115 0.515 31.445 0.845 ;
        RECT 31.12 -0.16 31.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.475 5.955 32.805 6.285 ;
        RECT 32.475 0.515 32.805 0.845 ;
        RECT 32.48 -0.16 32.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.835 5.955 34.165 6.285 ;
        RECT 33.835 0.515 34.165 0.845 ;
        RECT 33.84 -0.16 34.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.195 5.955 35.525 6.285 ;
        RECT 35.195 0.515 35.525 0.845 ;
        RECT 35.2 -0.16 35.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.555 5.955 36.885 6.285 ;
        RECT 36.555 0.515 36.885 0.845 ;
        RECT 36.56 -0.16 36.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.915 5.955 38.245 6.285 ;
        RECT 37.915 0.515 38.245 0.845 ;
        RECT 37.92 -0.16 38.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.275 5.955 39.605 6.285 ;
        RECT 39.275 0.515 39.605 0.845 ;
        RECT 39.28 -0.16 39.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.635 5.955 40.965 6.285 ;
        RECT 40.635 1.875 40.965 2.205 ;
        RECT 40.635 0.515 40.965 0.845 ;
        RECT 40.64 -0.16 40.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.995 5.955 42.325 6.285 ;
        RECT 41.995 1.875 42.325 2.205 ;
        RECT 41.995 0.515 42.325 0.845 ;
        RECT 42 -0.16 42.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.355 5.955 43.685 6.285 ;
        RECT 43.355 1.875 43.685 2.205 ;
        RECT 43.355 0.515 43.685 0.845 ;
        RECT 43.36 -0.16 43.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.715 5.955 45.045 6.285 ;
        RECT 44.715 0.515 45.045 0.845 ;
        RECT 44.72 -0.16 45.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.075 5.955 46.405 6.285 ;
        RECT 46.075 0.515 46.405 0.845 ;
        RECT 46.08 -0.16 46.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.435 5.955 47.765 6.285 ;
        RECT 47.435 0.515 47.765 0.845 ;
        RECT 47.44 -0.16 47.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.795 5.955 49.125 6.285 ;
        RECT 48.795 0.515 49.125 0.845 ;
        RECT 48.8 -0.16 49.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.155 5.955 50.485 6.285 ;
        RECT 50.155 0.515 50.485 0.845 ;
        RECT 50.16 -0.16 50.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.515 5.955 51.845 6.285 ;
        RECT 51.515 1.875 51.845 2.205 ;
        RECT 51.515 0.515 51.845 0.845 ;
        RECT 51.52 -0.16 51.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.875 5.955 53.205 6.285 ;
        RECT 52.875 1.875 53.205 2.205 ;
        RECT 52.875 0.515 53.205 0.845 ;
        RECT 52.88 -0.16 53.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.235 5.955 54.565 6.285 ;
        RECT 54.235 1.875 54.565 2.205 ;
        RECT 54.235 0.515 54.565 0.845 ;
        RECT 54.24 -0.16 54.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.595 5.955 55.925 6.285 ;
        RECT 55.595 0.515 55.925 0.845 ;
        RECT 55.6 -0.16 55.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.955 5.955 57.285 6.285 ;
        RECT 56.955 0.515 57.285 0.845 ;
        RECT 56.96 -0.16 57.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.315 5.955 58.645 6.285 ;
        RECT 58.315 0.515 58.645 0.845 ;
        RECT 58.32 -0.16 58.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.675 5.955 60.005 6.285 ;
        RECT 59.675 0.515 60.005 0.845 ;
        RECT 59.68 -0.16 60 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.035 5.955 61.365 6.285 ;
        RECT 61.035 0.515 61.365 0.845 ;
        RECT 61.04 -0.16 61.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.395 5.955 62.725 6.285 ;
        RECT 62.395 0.515 62.725 0.845 ;
        RECT 62.4 -0.16 62.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.755 5.955 64.085 6.285 ;
        RECT 63.755 1.875 64.085 2.205 ;
        RECT 63.755 0.515 64.085 0.845 ;
        RECT 63.76 -0.16 64.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.115 5.955 65.445 6.285 ;
        RECT 65.115 1.875 65.445 2.205 ;
        RECT 65.115 0.515 65.445 0.845 ;
        RECT 65.12 -0.16 65.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.475 5.955 66.805 6.285 ;
        RECT 66.475 1.875 66.805 2.205 ;
        RECT 66.475 0.515 66.805 0.845 ;
        RECT 66.48 -0.16 66.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.835 5.955 68.165 6.285 ;
        RECT 67.835 0.515 68.165 0.845 ;
        RECT 67.84 -0.16 68.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.195 5.955 69.525 6.285 ;
        RECT 69.195 0.515 69.525 0.845 ;
        RECT 69.2 -0.16 69.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.555 5.955 70.885 6.285 ;
        RECT 70.555 0.515 70.885 0.845 ;
        RECT 70.56 -0.16 70.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915 5.955 72.245 6.285 ;
        RECT 71.915 0.515 72.245 0.845 ;
        RECT 71.92 -0.16 72.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.275 5.955 73.605 6.285 ;
        RECT 73.275 0.515 73.605 0.845 ;
        RECT 73.28 -0.16 73.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.635 5.955 74.965 6.285 ;
        RECT 74.635 0.515 74.965 0.845 ;
        RECT 74.64 -0.16 74.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.995 5.955 76.325 6.285 ;
        RECT 75.995 1.875 76.325 2.205 ;
        RECT 75.995 0.515 76.325 0.845 ;
        RECT 76 -0.16 76.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.355 5.955 77.685 6.285 ;
        RECT 77.355 1.875 77.685 2.205 ;
        RECT 77.355 0.515 77.685 0.845 ;
        RECT 77.36 -0.16 77.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.715 5.955 79.045 6.285 ;
        RECT 78.715 1.875 79.045 2.205 ;
        RECT 78.715 0.515 79.045 0.845 ;
        RECT 78.72 -0.16 79.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.075 5.955 80.405 6.285 ;
        RECT 80.075 0.515 80.405 0.845 ;
        RECT 80.08 -0.16 80.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.435 5.955 81.765 6.285 ;
        RECT 81.435 0.515 81.765 0.845 ;
        RECT 81.44 -0.16 81.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.795 5.955 83.125 6.285 ;
        RECT 82.795 0.515 83.125 0.845 ;
        RECT 82.8 -0.16 83.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.155 5.955 84.485 6.285 ;
        RECT 84.155 0.515 84.485 0.845 ;
        RECT 84.16 -0.16 84.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.515 5.955 85.845 6.285 ;
        RECT 85.515 0.515 85.845 0.845 ;
        RECT 85.52 -0.16 85.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.875 5.955 87.205 6.285 ;
        RECT 86.875 0.515 87.205 0.845 ;
        RECT 86.88 -0.16 87.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.235 5.955 88.565 6.285 ;
        RECT 88.235 1.875 88.565 2.205 ;
        RECT 88.235 0.515 88.565 0.845 ;
        RECT 88.24 -0.16 88.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 89.595 5.955 89.925 6.285 ;
        RECT 89.595 1.875 89.925 2.205 ;
        RECT 89.595 0.515 89.925 0.845 ;
        RECT 89.6 -0.16 89.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.955 5.955 91.285 6.285 ;
        RECT 90.955 1.875 91.285 2.205 ;
        RECT 90.955 0.515 91.285 0.845 ;
        RECT 90.96 -0.16 91.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.315 5.955 92.645 6.285 ;
        RECT 92.315 0.515 92.645 0.845 ;
        RECT 92.32 -0.16 92.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.675 5.955 94.005 6.285 ;
        RECT 93.675 0.515 94.005 0.845 ;
        RECT 93.68 -0.16 94 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.035 5.955 95.365 6.285 ;
        RECT 95.035 0.515 95.365 0.845 ;
        RECT 95.04 -0.16 95.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.395 5.955 96.725 6.285 ;
        RECT 96.395 0.515 96.725 0.845 ;
        RECT 96.4 -0.16 96.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.755 5.955 98.085 6.285 ;
        RECT 97.755 0.515 98.085 0.845 ;
        RECT 97.76 -0.16 98.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.115 5.955 99.445 6.285 ;
        RECT 99.115 0.515 99.445 0.845 ;
        RECT 99.12 -0.16 99.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.475 5.955 100.805 6.285 ;
        RECT 100.475 1.875 100.805 2.205 ;
        RECT 100.475 0.515 100.805 0.845 ;
        RECT 100.48 -0.16 100.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.835 5.955 102.165 6.285 ;
        RECT 101.835 1.875 102.165 2.205 ;
        RECT 101.835 0.515 102.165 0.845 ;
        RECT 101.84 -0.16 102.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.195 5.955 103.525 6.285 ;
        RECT 103.195 1.875 103.525 2.205 ;
        RECT 103.195 0.515 103.525 0.845 ;
        RECT 103.2 -0.16 103.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 104.555 5.955 104.885 6.285 ;
        RECT 104.555 0.515 104.885 0.845 ;
        RECT 104.56 -0.16 104.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.915 5.955 106.245 6.285 ;
        RECT 105.915 0.515 106.245 0.845 ;
        RECT 105.92 -0.16 106.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.275 5.955 107.605 6.285 ;
        RECT 107.275 0.515 107.605 0.845 ;
        RECT 107.28 -0.16 107.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.635 5.955 108.965 6.285 ;
        RECT 108.635 0.515 108.965 0.845 ;
        RECT 108.64 -0.16 108.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.995 5.955 110.325 6.285 ;
        RECT 109.995 0.515 110.325 0.845 ;
        RECT 110 -0.16 110.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.355 5.955 111.685 6.285 ;
        RECT 111.355 0.515 111.685 0.845 ;
        RECT 111.36 -0.16 111.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.715 5.955 113.045 6.285 ;
        RECT 112.715 1.875 113.045 2.205 ;
        RECT 112.715 0.515 113.045 0.845 ;
        RECT 112.72 -0.16 113.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.075 5.955 114.405 6.285 ;
        RECT 114.075 1.875 114.405 2.205 ;
        RECT 114.075 0.515 114.405 0.845 ;
        RECT 114.08 -0.16 114.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.435 5.955 115.765 6.285 ;
        RECT 115.435 1.875 115.765 2.205 ;
        RECT 115.435 0.515 115.765 0.845 ;
        RECT 115.44 -0.16 115.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.795 5.955 117.125 6.285 ;
        RECT 116.795 0.515 117.125 0.845 ;
        RECT 116.8 -0.16 117.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.155 5.955 118.485 6.285 ;
        RECT 118.155 0.515 118.485 0.845 ;
        RECT 118.16 -0.16 118.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 119.515 5.955 119.845 6.285 ;
        RECT 119.515 0.515 119.845 0.845 ;
        RECT 119.52 -0.16 119.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.875 5.955 121.205 6.285 ;
        RECT 120.875 0.515 121.205 0.845 ;
        RECT 120.88 -0.16 121.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.235 5.955 122.565 6.285 ;
        RECT 122.235 0.515 122.565 0.845 ;
        RECT 122.24 -0.16 122.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.595 5.955 123.925 6.285 ;
        RECT 123.595 1.875 123.925 2.205 ;
        RECT 123.595 0.515 123.925 0.845 ;
        RECT 123.6 -0.16 123.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.955 5.955 125.285 6.285 ;
        RECT 124.955 1.875 125.285 2.205 ;
        RECT 124.955 0.515 125.285 0.845 ;
        RECT 124.96 -0.16 125.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.315 5.955 126.645 6.285 ;
        RECT 126.315 1.875 126.645 2.205 ;
        RECT 126.315 0.515 126.645 0.845 ;
        RECT 126.32 -0.16 126.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.675 5.955 128.005 6.285 ;
        RECT 127.675 0.515 128.005 0.845 ;
        RECT 127.68 -0.16 128 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.035 5.955 129.365 6.285 ;
        RECT 129.035 0.515 129.365 0.845 ;
        RECT 129.04 -0.16 129.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.395 5.955 130.725 6.285 ;
        RECT 130.395 0.515 130.725 0.845 ;
        RECT 130.4 -0.16 130.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.755 5.955 132.085 6.285 ;
        RECT 131.755 0.515 132.085 0.845 ;
        RECT 131.76 -0.16 132.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.115 5.955 133.445 6.285 ;
        RECT 133.115 0.515 133.445 0.845 ;
        RECT 133.12 -0.16 133.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.475 5.955 134.805 6.285 ;
        RECT 134.475 0.515 134.805 0.845 ;
        RECT 134.48 -0.16 134.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.835 5.955 136.165 6.285 ;
        RECT 135.835 1.875 136.165 2.205 ;
        RECT 135.835 0.515 136.165 0.845 ;
        RECT 135.84 -0.16 136.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.195 5.955 137.525 6.285 ;
        RECT 137.195 1.875 137.525 2.205 ;
        RECT 137.195 0.515 137.525 0.845 ;
        RECT 137.2 -0.16 137.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 138.555 5.955 138.885 6.285 ;
        RECT 138.555 1.875 138.885 2.205 ;
        RECT 138.555 0.515 138.885 0.845 ;
        RECT 138.56 -0.16 138.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.915 5.955 140.245 6.285 ;
        RECT 139.915 0.515 140.245 0.845 ;
        RECT 139.92 -0.16 140.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.275 5.955 141.605 6.285 ;
        RECT 141.275 0.515 141.605 0.845 ;
        RECT 141.28 -0.16 141.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.635 5.955 142.965 6.285 ;
        RECT 142.635 0.515 142.965 0.845 ;
        RECT 142.64 -0.16 142.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.995 5.955 144.325 6.285 ;
        RECT 143.995 0.515 144.325 0.845 ;
        RECT 144 -0.16 144.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.355 5.955 145.685 6.285 ;
        RECT 145.355 0.515 145.685 0.845 ;
        RECT 145.36 -0.16 145.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.715 5.955 147.045 6.285 ;
        RECT 146.715 0.515 147.045 0.845 ;
        RECT 146.72 -0.16 147.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.075 5.955 148.405 6.285 ;
        RECT 148.075 1.875 148.405 2.205 ;
        RECT 148.075 0.515 148.405 0.845 ;
        RECT 148.08 -0.16 148.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.435 5.955 149.765 6.285 ;
        RECT 149.435 1.875 149.765 2.205 ;
        RECT 149.435 0.515 149.765 0.845 ;
        RECT 149.44 -0.16 149.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.795 5.955 151.125 6.285 ;
        RECT 150.795 1.875 151.125 2.205 ;
        RECT 150.795 0.515 151.125 0.845 ;
        RECT 150.8 -0.16 151.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.155 5.955 152.485 6.285 ;
        RECT 152.155 0.515 152.485 0.845 ;
        RECT 152.16 -0.16 152.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.515 5.955 153.845 6.285 ;
        RECT 153.515 0.515 153.845 0.845 ;
        RECT 153.52 -0.16 153.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.875 5.955 155.205 6.285 ;
        RECT 154.875 0.515 155.205 0.845 ;
        RECT 154.88 -0.16 155.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.235 5.955 156.565 6.285 ;
        RECT 156.235 0.515 156.565 0.845 ;
        RECT 156.24 -0.16 156.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 157.595 5.955 157.925 6.285 ;
        RECT 157.595 0.515 157.925 0.845 ;
        RECT 157.6 -0.16 157.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.955 5.955 159.285 6.285 ;
        RECT 158.955 0.515 159.285 0.845 ;
        RECT 158.96 -0.16 159.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.315 5.955 160.645 6.285 ;
        RECT 160.315 1.875 160.645 2.205 ;
        RECT 160.315 0.515 160.645 0.845 ;
        RECT 160.32 -0.16 160.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.675 5.955 162.005 6.285 ;
        RECT 161.675 1.875 162.005 2.205 ;
        RECT 161.675 0.515 162.005 0.845 ;
        RECT 161.68 -0.16 162 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.035 5.955 163.365 6.285 ;
        RECT 163.035 1.875 163.365 2.205 ;
        RECT 163.035 0.515 163.365 0.845 ;
        RECT 163.04 -0.16 163.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 164.395 5.955 164.725 6.285 ;
        RECT 164.395 0.515 164.725 0.845 ;
        RECT 164.4 -0.16 164.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.755 5.955 166.085 6.285 ;
        RECT 165.755 0.515 166.085 0.845 ;
        RECT 165.76 -0.16 166.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.115 5.955 167.445 6.285 ;
        RECT 167.115 0.515 167.445 0.845 ;
        RECT 167.12 -0.16 167.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 168.475 5.955 168.805 6.285 ;
        RECT 168.475 0.515 168.805 0.845 ;
        RECT 168.48 -0.16 168.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.835 5.955 170.165 6.285 ;
        RECT 169.835 0.515 170.165 0.845 ;
        RECT 169.84 -0.16 170.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.195 5.955 171.525 6.285 ;
        RECT 171.195 0.515 171.525 0.845 ;
        RECT 171.2 -0.16 171.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.555 5.955 172.885 6.285 ;
        RECT 172.555 1.875 172.885 2.205 ;
        RECT 172.555 0.515 172.885 0.845 ;
        RECT 172.56 -0.16 172.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.915 5.955 174.245 6.285 ;
        RECT 173.915 1.875 174.245 2.205 ;
        RECT 173.915 0.515 174.245 0.845 ;
        RECT 173.92 -0.16 174.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.275 5.955 175.605 6.285 ;
        RECT 175.275 1.875 175.605 2.205 ;
        RECT 175.275 0.515 175.605 0.845 ;
        RECT 175.28 -0.16 175.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 176.635 5.955 176.965 6.285 ;
        RECT 176.635 0.515 176.965 0.845 ;
        RECT 176.64 -0.16 176.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.995 5.955 178.325 6.285 ;
        RECT 177.995 0.515 178.325 0.845 ;
        RECT 178 -0.16 178.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 179.355 5.955 179.685 6.285 ;
        RECT 179.355 0.515 179.685 0.845 ;
        RECT 179.36 -0.16 179.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.715 5.955 181.045 6.285 ;
        RECT 180.715 0.515 181.045 0.845 ;
        RECT 180.72 -0.16 181.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.075 5.955 182.405 6.285 ;
        RECT 182.075 0.515 182.405 0.845 ;
        RECT 182.08 -0.16 182.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 183.435 5.955 183.765 6.285 ;
        RECT 183.435 0.515 183.765 0.845 ;
        RECT 183.44 -0.16 183.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.795 5.955 185.125 6.285 ;
        RECT 184.795 1.875 185.125 2.205 ;
        RECT 184.795 0.515 185.125 0.845 ;
        RECT 184.8 -0.16 185.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.155 5.955 186.485 6.285 ;
        RECT 186.155 1.875 186.485 2.205 ;
        RECT 186.155 0.515 186.485 0.845 ;
        RECT 186.16 -0.16 186.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 187.515 5.955 187.845 6.285 ;
        RECT 187.515 1.875 187.845 2.205 ;
        RECT 187.515 0.515 187.845 0.845 ;
        RECT 187.52 -0.16 187.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.875 5.955 189.205 6.285 ;
        RECT 188.875 0.515 189.205 0.845 ;
        RECT 188.88 -0.16 189.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.235 5.955 190.565 6.285 ;
        RECT 190.235 0.515 190.565 0.845 ;
        RECT 190.24 -0.16 190.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 191.595 5.955 191.925 6.285 ;
        RECT 191.595 0.515 191.925 0.845 ;
        RECT 191.6 -0.16 191.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.955 5.955 193.285 6.285 ;
        RECT 192.955 0.515 193.285 0.845 ;
        RECT 192.96 -0.16 193.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.315 5.955 194.645 6.285 ;
        RECT 194.315 0.515 194.645 0.845 ;
        RECT 194.32 -0.16 194.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 195.675 5.955 196.005 6.285 ;
        RECT 195.675 1.875 196.005 2.205 ;
        RECT 195.675 0.515 196.005 0.845 ;
        RECT 195.68 -0.16 196 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.035 5.955 197.365 6.285 ;
        RECT 197.035 1.875 197.365 2.205 ;
        RECT 197.035 0.515 197.365 0.845 ;
        RECT 197.04 -0.16 197.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.395 5.955 198.725 6.285 ;
        RECT 198.395 1.875 198.725 2.205 ;
        RECT 198.395 0.515 198.725 0.845 ;
        RECT 198.4 -0.16 198.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.755 5.955 200.085 6.285 ;
        RECT 199.755 0.515 200.085 0.845 ;
        RECT 199.76 -0.16 200.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.115 5.955 201.445 6.285 ;
        RECT 201.115 0.515 201.445 0.845 ;
        RECT 201.12 -0.16 201.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 202.475 5.955 202.805 6.285 ;
        RECT 202.475 0.515 202.805 0.845 ;
        RECT 202.48 -0.16 202.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.835 5.955 204.165 6.285 ;
        RECT 203.835 0.515 204.165 0.845 ;
        RECT 203.84 -0.16 204.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.195 5.955 205.525 6.285 ;
        RECT 205.195 0.515 205.525 0.845 ;
        RECT 205.2 -0.16 205.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 206.555 5.955 206.885 6.285 ;
        RECT 206.555 0.515 206.885 0.845 ;
        RECT 206.56 -0.16 206.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.915 5.955 208.245 6.285 ;
        RECT 207.915 1.875 208.245 2.205 ;
        RECT 207.915 0.515 208.245 0.845 ;
        RECT 207.92 -0.16 208.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.275 5.955 209.605 6.285 ;
        RECT 209.275 1.875 209.605 2.205 ;
        RECT 209.275 0.515 209.605 0.845 ;
        RECT 209.28 -0.16 209.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 210.635 5.955 210.965 6.285 ;
        RECT 210.635 1.875 210.965 2.205 ;
        RECT 210.635 0.515 210.965 0.845 ;
        RECT 210.64 -0.16 210.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 211.995 5.955 212.325 6.285 ;
        RECT 211.995 0.515 212.325 0.845 ;
        RECT 212 -0.16 212.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 213.355 5.955 213.685 6.285 ;
        RECT 213.355 0.515 213.685 0.845 ;
        RECT 213.36 -0.16 213.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.715 5.955 215.045 6.285 ;
        RECT 214.715 0.515 215.045 0.845 ;
        RECT 214.72 -0.16 215.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.075 5.955 216.405 6.285 ;
        RECT 216.075 0.515 216.405 0.845 ;
        RECT 216.08 -0.16 216.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 217.435 5.955 217.765 6.285 ;
        RECT 217.435 0.515 217.765 0.845 ;
        RECT 217.44 -0.16 217.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.795 5.955 219.125 6.285 ;
        RECT 218.795 0.515 219.125 0.845 ;
        RECT 218.8 -0.16 219.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.155 5.955 220.485 6.285 ;
        RECT 220.155 1.875 220.485 2.205 ;
        RECT 220.155 0.515 220.485 0.845 ;
        RECT 220.16 -0.16 220.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 221.515 5.955 221.845 6.285 ;
        RECT 221.515 1.875 221.845 2.205 ;
        RECT 221.515 0.515 221.845 0.845 ;
        RECT 221.52 -0.16 221.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.875 5.955 223.205 6.285 ;
        RECT 222.875 1.875 223.205 2.205 ;
        RECT 222.875 0.515 223.205 0.845 ;
        RECT 222.88 -0.16 223.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 224.235 5.955 224.565 6.285 ;
        RECT 224.235 0.515 224.565 0.845 ;
        RECT 224.24 -0.16 224.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 225.595 5.955 225.925 6.285 ;
        RECT 225.595 0.515 225.925 0.845 ;
        RECT 225.6 -0.16 225.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.955 5.955 227.285 6.285 ;
        RECT 226.955 0.515 227.285 0.845 ;
        RECT 226.96 -0.16 227.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.315 5.955 228.645 6.285 ;
        RECT 228.315 0.515 228.645 0.845 ;
        RECT 228.32 -0.16 228.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 229.675 5.955 230.005 6.285 ;
        RECT 229.675 0.515 230.005 0.845 ;
        RECT 229.68 -0.16 230 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 231.035 5.955 231.365 6.285 ;
        RECT 231.035 0.515 231.365 0.845 ;
        RECT 231.04 -0.16 231.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 232.395 5.955 232.725 6.285 ;
        RECT 232.395 1.875 232.725 2.205 ;
        RECT 232.395 0.515 232.725 0.845 ;
        RECT 232.4 -0.16 232.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.755 5.955 234.085 6.285 ;
        RECT 233.755 1.875 234.085 2.205 ;
        RECT 233.755 0.515 234.085 0.845 ;
        RECT 233.76 -0.16 234.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 235.115 5.955 235.445 6.285 ;
        RECT 235.115 1.875 235.445 2.205 ;
        RECT 235.115 0.515 235.445 0.845 ;
        RECT 235.12 -0.16 235.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 236.475 5.955 236.805 6.285 ;
        RECT 236.475 0.515 236.805 0.845 ;
        RECT 236.48 -0.16 236.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 237.835 5.955 238.165 6.285 ;
        RECT 237.835 0.515 238.165 0.845 ;
        RECT 237.84 -0.16 238.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.195 5.955 239.525 6.285 ;
        RECT 239.195 0.515 239.525 0.845 ;
        RECT 239.2 -0.16 239.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 240.555 5.955 240.885 6.285 ;
        RECT 240.555 0.515 240.885 0.845 ;
        RECT 240.56 -0.16 240.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 241.915 5.955 242.245 6.285 ;
        RECT 241.915 0.515 242.245 0.845 ;
        RECT 241.92 -0.16 242.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 243.275 5.955 243.605 6.285 ;
        RECT 243.275 0.515 243.605 0.845 ;
        RECT 243.28 -0.16 243.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 244.635 5.955 244.965 6.285 ;
        RECT 244.635 1.875 244.965 2.205 ;
        RECT 244.635 0.515 244.965 0.845 ;
        RECT 244.64 -0.16 244.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 245.995 5.955 246.325 6.285 ;
        RECT 245.995 1.875 246.325 2.205 ;
        RECT 245.995 0.515 246.325 0.845 ;
        RECT 246 -0.16 246.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 247.355 5.955 247.685 6.285 ;
        RECT 247.355 1.875 247.685 2.205 ;
        RECT 247.355 0.515 247.685 0.845 ;
        RECT 247.36 -0.16 247.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.715 5.955 249.045 6.285 ;
        RECT 248.715 0.515 249.045 0.845 ;
        RECT 248.72 -0.16 249.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.075 5.955 250.405 6.285 ;
        RECT 250.075 0.515 250.405 0.845 ;
        RECT 250.08 -0.16 250.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 251.435 5.955 251.765 6.285 ;
        RECT 251.435 0.515 251.765 0.845 ;
        RECT 251.44 -0.16 251.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.795 5.955 253.125 6.285 ;
        RECT 252.795 0.515 253.125 0.845 ;
        RECT 252.8 -0.16 253.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 254.155 5.955 254.485 6.285 ;
        RECT 254.155 0.515 254.485 0.845 ;
        RECT 254.16 -0.16 254.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 255.515 5.955 255.845 6.285 ;
        RECT 255.515 1.875 255.845 2.205 ;
        RECT 255.515 0.515 255.845 0.845 ;
        RECT 255.52 -0.16 255.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 256.875 5.955 257.205 6.285 ;
        RECT 256.875 1.875 257.205 2.205 ;
        RECT 256.875 0.515 257.205 0.845 ;
        RECT 256.88 -0.16 257.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.235 5.955 258.565 6.285 ;
        RECT 258.235 1.875 258.565 2.205 ;
        RECT 258.235 0.515 258.565 0.845 ;
        RECT 258.24 -0.16 258.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 259.595 5.955 259.925 6.285 ;
        RECT 259.595 0.515 259.925 0.845 ;
        RECT 259.6 -0.16 259.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.955 5.955 261.285 6.285 ;
        RECT 260.955 0.515 261.285 0.845 ;
        RECT 260.96 -0.16 261.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.315 5.955 262.645 6.285 ;
        RECT 262.315 0.515 262.645 0.845 ;
        RECT 262.32 -0.16 262.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 263.675 5.955 264.005 6.285 ;
        RECT 263.675 0.515 264.005 0.845 ;
        RECT 263.68 -0.16 264 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 265.035 5.955 265.365 6.285 ;
        RECT 265.035 0.515 265.365 0.845 ;
        RECT 265.04 -0.16 265.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 266.395 5.955 266.725 6.285 ;
        RECT 266.395 0.515 266.725 0.845 ;
        RECT 266.4 -0.16 266.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 267.755 5.955 268.085 6.285 ;
        RECT 267.755 1.875 268.085 2.205 ;
        RECT 267.755 0.515 268.085 0.845 ;
        RECT 267.76 -0.16 268.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.115 5.955 269.445 6.285 ;
        RECT 269.115 1.875 269.445 2.205 ;
        RECT 269.115 0.515 269.445 0.845 ;
        RECT 269.12 -0.16 269.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 270.475 5.955 270.805 6.285 ;
        RECT 270.475 1.875 270.805 2.205 ;
        RECT 270.475 0.515 270.805 0.845 ;
        RECT 270.48 -0.16 270.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.835 5.955 272.165 6.285 ;
        RECT 271.835 0.515 272.165 0.845 ;
        RECT 271.84 -0.16 272.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.195 5.955 273.525 6.285 ;
        RECT 273.195 0.515 273.525 0.845 ;
        RECT 273.2 -0.16 273.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 274.555 5.955 274.885 6.285 ;
        RECT 274.555 0.515 274.885 0.845 ;
        RECT 274.56 -0.16 274.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.915 5.955 276.245 6.285 ;
        RECT 275.915 0.515 276.245 0.845 ;
        RECT 275.92 -0.16 276.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 277.275 5.955 277.605 6.285 ;
        RECT 277.275 0.515 277.605 0.845 ;
        RECT 277.28 -0.16 277.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 278.635 5.955 278.965 6.285 ;
        RECT 278.635 0.515 278.965 0.845 ;
        RECT 278.64 -0.16 278.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.995 5.955 280.325 6.285 ;
        RECT 279.995 1.875 280.325 2.205 ;
        RECT 279.995 0.515 280.325 0.845 ;
        RECT 280 -0.16 280.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 281.355 5.955 281.685 6.285 ;
        RECT 281.355 1.875 281.685 2.205 ;
        RECT 281.355 0.515 281.685 0.845 ;
        RECT 281.36 -0.16 281.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.715 5.955 283.045 6.285 ;
        RECT 282.715 1.875 283.045 2.205 ;
        RECT 282.715 0.515 283.045 0.845 ;
        RECT 282.72 -0.16 283.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 284.075 5.955 284.405 6.285 ;
        RECT 284.075 0.515 284.405 0.845 ;
        RECT 284.08 -0.16 284.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 285.435 5.955 285.765 6.285 ;
        RECT 285.435 0.515 285.765 0.845 ;
        RECT 285.44 -0.16 285.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.795 5.955 287.125 6.285 ;
        RECT 286.795 0.515 287.125 0.845 ;
        RECT 286.8 -0.16 287.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.155 5.955 288.485 6.285 ;
        RECT 288.155 0.515 288.485 0.845 ;
        RECT 288.16 -0.16 288.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 289.515 5.955 289.845 6.285 ;
        RECT 289.515 0.515 289.845 0.845 ;
        RECT 289.52 -0.16 289.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.875 5.955 291.205 6.285 ;
        RECT 290.875 0.515 291.205 0.845 ;
        RECT 290.88 -0.16 291.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.235 5.955 292.565 6.285 ;
        RECT 292.235 1.875 292.565 2.205 ;
        RECT 292.235 0.515 292.565 0.845 ;
        RECT 292.24 -0.16 292.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 293.595 5.955 293.925 6.285 ;
        RECT 293.595 1.875 293.925 2.205 ;
        RECT 293.595 0.515 293.925 0.845 ;
        RECT 293.6 -0.16 293.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.955 5.955 295.285 6.285 ;
        RECT 294.955 1.875 295.285 2.205 ;
        RECT 294.955 0.515 295.285 0.845 ;
        RECT 294.96 -0.16 295.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 296.315 5.955 296.645 6.285 ;
        RECT 296.315 0.515 296.645 0.845 ;
        RECT 296.32 -0.16 296.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 297.675 5.955 298.005 6.285 ;
        RECT 297.675 0.515 298.005 0.845 ;
        RECT 297.68 -0.16 298 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 299.035 5.955 299.365 6.285 ;
        RECT 299.035 0.515 299.365 0.845 ;
        RECT 299.04 -0.16 299.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 300.395 5.955 300.725 6.285 ;
        RECT 300.395 0.515 300.725 0.845 ;
        RECT 300.4 -0.16 300.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.755 5.955 302.085 6.285 ;
        RECT 301.755 0.515 302.085 0.845 ;
        RECT 301.76 -0.16 302.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.115 5.955 303.445 6.285 ;
        RECT 303.115 0.515 303.445 0.845 ;
        RECT 303.12 -0.16 303.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 304.475 5.955 304.805 6.285 ;
        RECT 304.475 1.875 304.805 2.205 ;
        RECT 304.475 0.515 304.805 0.845 ;
        RECT 304.48 -0.16 304.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.835 5.955 306.165 6.285 ;
        RECT 305.835 1.875 306.165 2.205 ;
        RECT 305.835 0.515 306.165 0.845 ;
        RECT 305.84 -0.16 306.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.195 5.955 307.525 6.285 ;
        RECT 307.195 1.875 307.525 2.205 ;
        RECT 307.195 0.515 307.525 0.845 ;
        RECT 307.2 -0.16 307.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 308.555 5.955 308.885 6.285 ;
        RECT 308.555 0.515 308.885 0.845 ;
        RECT 308.56 -0.16 308.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.915 5.955 310.245 6.285 ;
        RECT 309.915 0.515 310.245 0.845 ;
        RECT 309.92 -0.16 310.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 311.275 5.955 311.605 6.285 ;
        RECT 311.275 0.515 311.605 0.845 ;
        RECT 311.28 -0.16 311.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 312.635 5.955 312.965 6.285 ;
        RECT 312.635 0.515 312.965 0.845 ;
        RECT 312.64 -0.16 312.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.995 5.955 314.325 6.285 ;
        RECT 313.995 0.515 314.325 0.845 ;
        RECT 314 -0.16 314.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 315.355 5.955 315.685 6.285 ;
        RECT 315.355 0.515 315.685 0.845 ;
        RECT 315.36 -0.16 315.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 316.715 5.955 317.045 6.285 ;
        RECT 316.715 1.875 317.045 2.205 ;
        RECT 316.715 0.515 317.045 0.845 ;
        RECT 316.72 -0.16 317.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.075 5.955 318.405 6.285 ;
        RECT 318.075 1.875 318.405 2.205 ;
        RECT 318.075 0.515 318.405 0.845 ;
        RECT 318.08 -0.16 318.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 319.435 5.955 319.765 6.285 ;
        RECT 319.435 1.875 319.765 2.205 ;
        RECT 319.435 0.515 319.765 0.845 ;
        RECT 319.44 -0.16 319.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 320.795 5.955 321.125 6.285 ;
        RECT 320.795 0.515 321.125 0.845 ;
        RECT 320.8 -0.16 321.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 322.155 5.955 322.485 6.285 ;
        RECT 322.155 0.515 322.485 0.845 ;
        RECT 322.16 -0.16 322.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 323.515 5.955 323.845 6.285 ;
        RECT 323.515 0.515 323.845 0.845 ;
        RECT 323.52 -0.16 323.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.875 5.955 325.205 6.285 ;
        RECT 324.875 0.515 325.205 0.845 ;
        RECT 324.88 -0.16 325.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 326.235 5.955 326.565 6.285 ;
        RECT 326.235 0.515 326.565 0.845 ;
        RECT 326.24 -0.16 326.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 327.595 5.955 327.925 6.285 ;
        RECT 327.595 1.875 327.925 2.205 ;
        RECT 327.595 0.515 327.925 0.845 ;
        RECT 327.6 -0.16 327.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 328.955 5.955 329.285 6.285 ;
        RECT 328.955 1.875 329.285 2.205 ;
        RECT 328.955 0.515 329.285 0.845 ;
        RECT 328.96 -0.16 329.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.315 5.955 330.645 6.285 ;
        RECT 330.315 1.875 330.645 2.205 ;
        RECT 330.315 0.515 330.645 0.845 ;
        RECT 330.32 -0.16 330.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 331.675 5.955 332.005 6.285 ;
        RECT 331.675 0.515 332.005 0.845 ;
        RECT 331.68 -0.16 332 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 333.035 5.955 333.365 6.285 ;
        RECT 333.035 0.515 333.365 0.845 ;
        RECT 333.04 -0.16 333.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 334.395 5.955 334.725 6.285 ;
        RECT 334.395 0.515 334.725 0.845 ;
        RECT 334.4 -0.16 334.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.755 5.955 336.085 6.285 ;
        RECT 335.755 0.515 336.085 0.845 ;
        RECT 335.76 -0.16 336.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 337.115 5.955 337.445 6.285 ;
        RECT 337.115 0.515 337.445 0.845 ;
        RECT 337.12 -0.16 337.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 338.475 5.955 338.805 6.285 ;
        RECT 338.475 0.515 338.805 0.845 ;
        RECT 338.48 -0.16 338.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 339.835 5.955 340.165 6.285 ;
        RECT 339.835 1.875 340.165 2.205 ;
        RECT 339.835 0.515 340.165 0.845 ;
        RECT 339.84 -0.16 340.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 341.195 5.955 341.525 6.285 ;
        RECT 341.195 1.875 341.525 2.205 ;
        RECT 341.195 0.515 341.525 0.845 ;
        RECT 341.2 -0.16 341.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 342.555 5.955 342.885 6.285 ;
        RECT 342.555 1.875 342.885 2.205 ;
        RECT 342.555 0.515 342.885 0.845 ;
        RECT 342.56 -0.16 342.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 343.915 5.955 344.245 6.285 ;
        RECT 343.915 0.515 344.245 0.845 ;
        RECT 343.92 -0.16 344.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 345.275 5.955 345.605 6.285 ;
        RECT 345.275 0.515 345.605 0.845 ;
        RECT 345.28 -0.16 345.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 346.635 5.955 346.965 6.285 ;
        RECT 346.635 0.515 346.965 0.845 ;
        RECT 346.64 -0.16 346.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 347.995 5.955 348.325 6.285 ;
        RECT 347.995 0.515 348.325 0.845 ;
        RECT 348 -0.16 348.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 349.355 5.955 349.685 6.285 ;
        RECT 349.355 0.515 349.685 0.845 ;
        RECT 349.36 -0.16 349.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 350.715 5.955 351.045 6.285 ;
        RECT 350.715 0.515 351.045 0.845 ;
        RECT 350.72 -0.16 351.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 352.075 5.955 352.405 6.285 ;
        RECT 352.075 1.875 352.405 2.205 ;
        RECT 352.075 0.515 352.405 0.845 ;
        RECT 352.08 -0.16 352.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 353.435 5.955 353.765 6.285 ;
        RECT 353.435 1.875 353.765 2.205 ;
        RECT 353.435 0.515 353.765 0.845 ;
        RECT 353.44 -0.16 353.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.795 5.955 355.125 6.285 ;
        RECT 354.795 1.875 355.125 2.205 ;
        RECT 354.795 0.515 355.125 0.845 ;
        RECT 354.8 -0.16 355.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 356.155 5.955 356.485 6.285 ;
        RECT 356.155 0.515 356.485 0.845 ;
        RECT 356.16 -0.16 356.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 357.515 5.955 357.845 6.285 ;
        RECT 357.515 0.515 357.845 0.845 ;
        RECT 357.52 -0.16 357.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 358.875 5.955 359.205 6.285 ;
        RECT 358.875 0.515 359.205 0.845 ;
        RECT 358.88 -0.16 359.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 360.235 5.955 360.565 6.285 ;
        RECT 360.235 0.515 360.565 0.845 ;
        RECT 360.24 -0.16 360.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 361.595 5.955 361.925 6.285 ;
        RECT 361.595 0.515 361.925 0.845 ;
        RECT 361.6 -0.16 361.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 362.955 5.955 363.285 6.285 ;
        RECT 362.955 0.515 363.285 0.845 ;
        RECT 362.96 -0.16 363.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 364.315 5.955 364.645 6.285 ;
        RECT 364.315 1.875 364.645 2.205 ;
        RECT 364.315 0.515 364.645 0.845 ;
        RECT 364.32 -0.16 364.64 7.64 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 321.475 1.195 321.805 1.525 ;
        RECT 321.475 -0.165 321.805 0.165 ;
        RECT 321.48 -0.165 321.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 322.835 1.195 323.165 1.525 ;
        RECT 322.835 -0.165 323.165 0.165 ;
        RECT 322.84 -0.165 323.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.195 1.195 324.525 1.525 ;
        RECT 324.195 -0.165 324.525 0.165 ;
        RECT 324.2 -0.165 324.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 325.555 1.195 325.885 1.525 ;
        RECT 325.555 -0.165 325.885 0.165 ;
        RECT 325.56 -0.165 325.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 326.915 1.195 327.245 1.525 ;
        RECT 326.915 -0.165 327.245 0.165 ;
        RECT 326.92 -0.165 327.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 328.275 1.195 328.605 1.525 ;
        RECT 328.275 -0.165 328.605 0.165 ;
        RECT 328.28 -0.165 328.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 329.635 1.195 329.965 1.525 ;
        RECT 329.635 -0.165 329.965 0.165 ;
        RECT 329.64 -0.165 329.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.995 1.195 331.325 1.525 ;
        RECT 330.995 -0.165 331.325 0.165 ;
        RECT 331 -0.165 331.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 332.355 1.195 332.685 1.525 ;
        RECT 332.355 -0.165 332.685 0.165 ;
        RECT 332.36 -0.165 332.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 333.715 1.195 334.045 1.525 ;
        RECT 333.715 -0.165 334.045 0.165 ;
        RECT 333.72 -0.165 334.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.075 1.195 335.405 1.525 ;
        RECT 335.075 -0.165 335.405 0.165 ;
        RECT 335.08 -0.165 335.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 336.435 1.195 336.765 1.525 ;
        RECT 336.435 -0.165 336.765 0.165 ;
        RECT 336.44 -0.165 336.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 337.795 1.195 338.125 1.525 ;
        RECT 337.795 -0.165 338.125 0.165 ;
        RECT 337.8 -0.165 338.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 339.155 1.195 339.485 1.525 ;
        RECT 339.155 -0.165 339.485 0.165 ;
        RECT 339.16 -0.165 339.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 340.515 1.195 340.845 1.525 ;
        RECT 340.515 -0.165 340.845 0.165 ;
        RECT 340.52 -0.165 340.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 341.875 1.195 342.205 1.525 ;
        RECT 341.875 -0.165 342.205 0.165 ;
        RECT 341.88 -0.165 342.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 343.235 1.195 343.565 1.525 ;
        RECT 343.235 -0.165 343.565 0.165 ;
        RECT 343.24 -0.165 343.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 344.595 1.195 344.925 1.525 ;
        RECT 344.595 -0.165 344.925 0.165 ;
        RECT 344.6 -0.165 344.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 345.955 1.195 346.285 1.525 ;
        RECT 345.955 -0.165 346.285 0.165 ;
        RECT 345.96 -0.165 346.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 347.315 1.195 347.645 1.525 ;
        RECT 347.315 -0.165 347.645 0.165 ;
        RECT 347.32 -0.165 347.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 348.675 1.195 349.005 1.525 ;
        RECT 348.675 -0.165 349.005 0.165 ;
        RECT 348.68 -0.165 349 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 350.035 1.195 350.365 1.525 ;
        RECT 350.035 -0.165 350.365 0.165 ;
        RECT 350.04 -0.165 350.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 351.395 1.195 351.725 1.525 ;
        RECT 351.395 -0.165 351.725 0.165 ;
        RECT 351.4 -0.165 351.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 352.755 1.195 353.085 1.525 ;
        RECT 352.755 -0.165 353.085 0.165 ;
        RECT 352.76 -0.165 353.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.115 1.195 354.445 1.525 ;
        RECT 354.115 -0.165 354.445 0.165 ;
        RECT 354.12 -0.165 354.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 355.475 1.195 355.805 1.525 ;
        RECT 355.475 -0.165 355.805 0.165 ;
        RECT 355.48 -0.165 355.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 356.835 1.195 357.165 1.525 ;
        RECT 356.835 -0.165 357.165 0.165 ;
        RECT 356.84 -0.165 357.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 358.195 1.195 358.525 1.525 ;
        RECT 358.195 -0.165 358.525 0.165 ;
        RECT 358.2 -0.165 358.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 359.555 1.195 359.885 1.525 ;
        RECT 359.555 -0.165 359.885 0.165 ;
        RECT 359.56 -0.165 359.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 360.915 1.195 361.245 1.525 ;
        RECT 360.915 -0.165 361.245 0.165 ;
        RECT 360.92 -0.165 361.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 362.275 1.195 362.605 1.525 ;
        RECT 362.275 -0.165 362.605 0.165 ;
        RECT 362.28 -0.165 362.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 363.635 1.195 363.965 1.525 ;
        RECT 363.635 -0.165 363.965 0.165 ;
        RECT 363.64 -0.165 363.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 364.995 1.195 365.325 1.525 ;
        RECT 364.995 -0.165 365.325 0.165 ;
        RECT 365 -0.165 365.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 366.355 1.195 366.685 1.525 ;
        RECT 366.355 -0.165 366.685 0.165 ;
        RECT 366.36 -0.165 366.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 367.715 1.195 368.045 1.525 ;
        RECT 367.715 -0.165 368.045 0.165 ;
        RECT 367.72 -0.165 368.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 369.075 1.195 369.405 1.525 ;
        RECT 369.075 -0.165 369.405 0.165 ;
        RECT 369.08 -0.165 369.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 370.435 1.195 370.765 1.525 ;
        RECT 370.435 -0.165 370.765 0.165 ;
        RECT 370.44 -0.165 370.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 371.795 1.195 372.125 1.525 ;
        RECT 371.795 -0.165 372.125 0.165 ;
        RECT 371.8 -0.165 372.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 373.155 1.195 373.485 1.525 ;
        RECT 373.155 -0.165 373.485 0.165 ;
        RECT 373.16 -0.165 373.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 374.515 1.195 374.845 1.525 ;
        RECT 374.515 -0.165 374.845 0.165 ;
        RECT 374.52 -0.165 374.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 375.875 1.195 376.205 1.525 ;
        RECT 375.875 -0.165 376.205 0.165 ;
        RECT 375.88 -0.165 376.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 377.235 1.195 377.565 1.525 ;
        RECT 377.235 -0.165 377.565 0.165 ;
        RECT 377.24 -0.165 377.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 378.595 1.195 378.925 1.525 ;
        RECT 378.595 -0.165 378.925 0.165 ;
        RECT 378.6 -0.165 378.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 379.955 1.195 380.285 1.525 ;
        RECT 379.955 -0.165 380.285 0.165 ;
        RECT 379.96 -0.165 380.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 381.315 1.195 381.645 1.525 ;
        RECT 381.315 -0.165 381.645 0.165 ;
        RECT 381.32 -0.165 381.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 382.675 1.195 383.005 1.525 ;
        RECT 382.675 -0.165 383.005 0.165 ;
        RECT 382.68 -0.165 383 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 384.035 1.195 384.365 1.525 ;
        RECT 384.035 -0.165 384.365 0.165 ;
        RECT 384.04 -0.165 384.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 385.395 1.195 385.725 1.525 ;
        RECT 385.395 -0.165 385.725 0.165 ;
        RECT 385.4 -0.165 385.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 386.755 1.195 387.085 1.525 ;
        RECT 386.755 -0.165 387.085 0.165 ;
        RECT 386.76 -0.165 387.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 388.115 1.195 388.445 1.525 ;
        RECT 388.115 -0.165 388.445 0.165 ;
        RECT 388.12 -0.165 388.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 389.475 1.195 389.805 1.525 ;
        RECT 389.475 -0.165 389.805 0.165 ;
        RECT 389.48 -0.165 389.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 390.835 1.195 391.165 1.525 ;
        RECT 390.835 -0.165 391.165 0.165 ;
        RECT 390.84 -0.165 391.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 392.195 1.195 392.525 1.525 ;
        RECT 392.195 -0.165 392.525 0.165 ;
        RECT 392.2 -0.165 392.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 393.555 1.195 393.885 1.525 ;
        RECT 393.555 -0.165 393.885 0.165 ;
        RECT 393.56 -0.165 393.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 394.915 1.195 395.245 1.525 ;
        RECT 394.915 -0.165 395.245 0.165 ;
        RECT 394.92 -0.165 395.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 396.275 1.195 396.605 1.525 ;
        RECT 396.275 -0.165 396.605 0.165 ;
        RECT 396.28 -0.165 396.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 397.635 1.195 397.965 1.525 ;
        RECT 397.635 -0.165 397.965 0.165 ;
        RECT 397.64 -0.165 397.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 398.995 1.195 399.325 1.525 ;
        RECT 398.995 -0.165 399.325 0.165 ;
        RECT 399 -0.165 399.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 400.355 1.195 400.685 1.525 ;
        RECT 400.355 -0.165 400.685 0.165 ;
        RECT 400.36 -0.165 400.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 401.715 1.195 402.045 1.525 ;
        RECT 401.715 -0.165 402.045 0.165 ;
        RECT 401.72 -0.165 402.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 403.075 1.195 403.405 1.525 ;
        RECT 403.075 -0.165 403.405 0.165 ;
        RECT 403.08 -0.165 403.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 404.435 1.195 404.765 1.525 ;
        RECT 404.435 -0.165 404.765 0.165 ;
        RECT 404.44 -0.165 404.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 405.795 1.195 406.125 1.525 ;
        RECT 405.795 -0.165 406.125 0.165 ;
        RECT 405.8 -0.165 406.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 407.155 1.195 407.485 1.525 ;
        RECT 407.155 -0.165 407.485 0.165 ;
        RECT 407.16 -0.165 407.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 408.515 1.195 408.845 1.525 ;
        RECT 408.515 -0.165 408.845 0.165 ;
        RECT 408.52 -0.165 408.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 409.875 1.195 410.205 1.525 ;
        RECT 409.875 -0.165 410.205 0.165 ;
        RECT 409.88 -0.165 410.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 411.235 1.195 411.565 1.525 ;
        RECT 411.235 -0.165 411.565 0.165 ;
        RECT 411.24 -0.165 411.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 412.595 1.195 412.925 1.525 ;
        RECT 412.595 -0.165 412.925 0.165 ;
        RECT 412.6 -0.165 412.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 413.955 1.195 414.285 1.525 ;
        RECT 413.955 -0.165 414.285 0.165 ;
        RECT 413.96 -0.165 414.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 415.315 1.195 415.645 1.525 ;
        RECT 415.315 -0.165 415.645 0.165 ;
        RECT 415.32 -0.165 415.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 416.675 1.195 417.005 1.525 ;
        RECT 416.675 -0.165 417.005 0.165 ;
        RECT 416.68 -0.165 417 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 418.035 1.195 418.365 1.525 ;
        RECT 418.035 -0.165 418.365 0.165 ;
        RECT 418.04 -0.165 418.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 419.395 1.195 419.725 1.525 ;
        RECT 419.395 -0.165 419.725 0.165 ;
        RECT 419.4 -0.165 419.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 420.755 1.195 421.085 1.525 ;
        RECT 420.755 -0.165 421.085 0.165 ;
        RECT 420.76 -0.165 421.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 422.115 1.195 422.445 1.525 ;
        RECT 422.115 -0.165 422.445 0.165 ;
        RECT 422.12 -0.165 422.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 423.475 1.195 423.805 1.525 ;
        RECT 423.475 -0.165 423.805 0.165 ;
        RECT 423.48 -0.165 423.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 424.835 1.195 425.165 1.525 ;
        RECT 424.835 -0.165 425.165 0.165 ;
        RECT 424.84 -0.165 425.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 426.195 1.195 426.525 1.525 ;
        RECT 426.195 -0.165 426.525 0.165 ;
        RECT 426.2 -0.165 426.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 427.555 1.195 427.885 1.525 ;
        RECT 427.555 -0.165 427.885 0.165 ;
        RECT 427.56 -0.165 427.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 428.915 1.195 429.245 1.525 ;
        RECT 428.915 -0.165 429.245 0.165 ;
        RECT 428.92 -0.165 429.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 430.275 1.195 430.605 1.525 ;
        RECT 430.275 -0.165 430.605 0.165 ;
        RECT 430.28 -0.165 430.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 431.635 1.195 431.965 1.525 ;
        RECT 431.635 -0.165 431.965 0.165 ;
        RECT 431.64 -0.165 431.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 432.995 1.195 433.325 1.525 ;
        RECT 432.995 -0.165 433.325 0.165 ;
        RECT 433 -0.165 433.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 434.355 1.195 434.685 1.525 ;
        RECT 434.355 -0.165 434.685 0.165 ;
        RECT 434.36 -0.165 434.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 435.715 1.195 436.045 1.525 ;
        RECT 435.715 -0.165 436.045 0.165 ;
        RECT 435.72 -0.165 436.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 437.075 1.195 437.405 1.525 ;
        RECT 437.075 -0.165 437.405 0.165 ;
        RECT 437.08 -0.165 437.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 438.435 1.195 438.765 1.525 ;
        RECT 438.435 -0.165 438.765 0.165 ;
        RECT 438.44 -0.165 438.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 439.795 1.195 440.125 1.525 ;
        RECT 439.795 -0.165 440.125 0.165 ;
        RECT 439.8 -0.165 440.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 441.155 1.195 441.485 1.525 ;
        RECT 441.155 -0.165 441.485 0.165 ;
        RECT 441.16 -0.165 441.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 442.515 1.195 442.845 1.525 ;
        RECT 442.515 -0.165 442.845 0.165 ;
        RECT 442.52 -0.165 442.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 443.875 1.195 444.205 1.525 ;
        RECT 443.875 -0.165 444.205 0.165 ;
        RECT 443.88 -0.165 444.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 445.235 1.195 445.565 1.525 ;
        RECT 445.235 -0.165 445.565 0.165 ;
        RECT 445.24 -0.165 445.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 446.595 1.195 446.925 1.525 ;
        RECT 446.595 -0.165 446.925 0.165 ;
        RECT 446.6 -0.165 446.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 447.955 1.195 448.285 1.525 ;
        RECT 447.955 -0.165 448.285 0.165 ;
        RECT 447.96 -0.165 448.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 449.315 1.195 449.645 1.525 ;
        RECT 449.315 -0.165 449.645 0.165 ;
        RECT 449.32 -0.165 449.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 450.675 1.195 451.005 1.525 ;
        RECT 450.675 -0.165 451.005 0.165 ;
        RECT 450.68 -0.165 451 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 452.035 1.195 452.365 1.525 ;
        RECT 452.035 -0.165 452.365 0.165 ;
        RECT 452.04 -0.165 452.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 453.395 1.195 453.725 1.525 ;
        RECT 453.395 -0.165 453.725 0.165 ;
        RECT 453.4 -0.165 453.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 454.755 1.195 455.085 1.525 ;
        RECT 454.755 -0.165 455.085 0.165 ;
        RECT 454.76 -0.165 455.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 456.115 1.195 456.445 1.525 ;
        RECT 456.115 -0.165 456.445 0.165 ;
        RECT 456.12 -0.165 456.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 457.475 1.195 457.805 1.525 ;
        RECT 457.475 -0.165 457.805 0.165 ;
        RECT 457.48 -0.165 457.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 458.835 1.195 459.165 1.525 ;
        RECT 458.835 -0.165 459.165 0.165 ;
        RECT 458.84 -0.165 459.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 460.195 1.195 460.525 1.525 ;
        RECT 460.195 -0.165 460.525 0.165 ;
        RECT 460.2 -0.165 460.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 461.555 1.195 461.885 1.525 ;
        RECT 461.555 -0.165 461.885 0.165 ;
        RECT 461.56 -0.165 461.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 462.915 1.195 463.245 1.525 ;
        RECT 462.915 -0.165 463.245 0.165 ;
        RECT 462.92 -0.165 463.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 464.275 1.195 464.605 1.525 ;
        RECT 464.275 -0.165 464.605 0.165 ;
        RECT 464.28 -0.165 464.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 465.635 1.195 465.965 1.525 ;
        RECT 465.635 -0.165 465.965 0.165 ;
        RECT 465.64 -0.165 465.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 466.995 1.195 467.325 1.525 ;
        RECT 466.995 -0.165 467.325 0.165 ;
        RECT 467 -0.165 467.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 468.355 1.195 468.685 1.525 ;
        RECT 468.355 -0.165 468.685 0.165 ;
        RECT 468.36 -0.165 468.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 469.715 1.195 470.045 1.525 ;
        RECT 469.715 -0.165 470.045 0.165 ;
        RECT 469.72 -0.165 470.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 471.075 1.195 471.405 1.525 ;
        RECT 471.075 -0.165 471.405 0.165 ;
        RECT 471.08 -0.165 471.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 472.435 1.195 472.765 1.525 ;
        RECT 472.435 -0.165 472.765 0.165 ;
        RECT 472.44 -0.165 472.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 473.795 1.195 474.125 1.525 ;
        RECT 473.795 -0.165 474.125 0.165 ;
        RECT 473.8 -0.165 474.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 475.155 1.195 475.485 1.525 ;
        RECT 475.155 -0.165 475.485 0.165 ;
        RECT 475.16 -0.165 475.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 476.515 1.195 476.845 1.525 ;
        RECT 476.515 -0.165 476.845 0.165 ;
        RECT 476.52 -0.165 476.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 477.875 1.195 478.205 1.525 ;
        RECT 477.875 -0.165 478.205 0.165 ;
        RECT 477.88 -0.165 478.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 479.235 1.195 479.565 1.525 ;
        RECT 479.235 -0.165 479.565 0.165 ;
        RECT 479.24 -0.165 479.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 480.595 1.195 480.925 1.525 ;
        RECT 480.595 -0.165 480.925 0.165 ;
        RECT 480.6 -0.165 480.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 481.955 1.195 482.285 1.525 ;
        RECT 481.955 -0.165 482.285 0.165 ;
        RECT 481.96 -0.165 482.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 483.315 1.195 483.645 1.525 ;
        RECT 483.315 -0.165 483.645 0.165 ;
        RECT 483.32 -0.165 483.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 484.675 1.195 485.005 1.525 ;
        RECT 484.675 -0.165 485.005 0.165 ;
        RECT 484.68 -0.165 485 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 486.035 1.195 486.365 1.525 ;
        RECT 486.035 -0.165 486.365 0.165 ;
        RECT 486.04 -0.165 486.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 487.395 1.195 487.725 1.525 ;
        RECT 487.395 -0.165 487.725 0.165 ;
        RECT 487.4 -0.165 487.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 488.755 1.195 489.085 1.525 ;
        RECT 488.755 -0.165 489.085 0.165 ;
        RECT 488.76 -0.165 489.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 490.115 1.195 490.445 1.525 ;
        RECT 490.115 -0.165 490.445 0.165 ;
        RECT 490.12 -0.165 490.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 491.475 1.195 491.805 1.525 ;
        RECT 491.475 -0.165 491.805 0.165 ;
        RECT 491.48 -0.165 491.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 492.835 1.195 493.165 1.525 ;
        RECT 492.835 -0.165 493.165 0.165 ;
        RECT 492.84 -0.165 493.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 494.195 1.195 494.525 1.525 ;
        RECT 494.195 -0.165 494.525 0.165 ;
        RECT 494.2 -0.165 494.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 495.555 1.195 495.885 1.525 ;
        RECT 495.555 -0.165 495.885 0.165 ;
        RECT 495.56 -0.165 495.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 496.915 1.195 497.245 1.525 ;
        RECT 496.915 -0.165 497.245 0.165 ;
        RECT 496.92 -0.165 497.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 498.275 1.195 498.605 1.525 ;
        RECT 498.275 -0.165 498.605 0.165 ;
        RECT 498.28 -0.165 498.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 499.635 1.195 499.965 1.525 ;
        RECT 499.635 -0.165 499.965 0.165 ;
        RECT 499.64 -0.165 499.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 500.995 1.195 501.325 1.525 ;
        RECT 500.995 -0.165 501.325 0.165 ;
        RECT 501 -0.165 501.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 502.355 1.195 502.685 1.525 ;
        RECT 502.355 -0.165 502.685 0.165 ;
        RECT 502.36 -0.165 502.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 503.715 1.195 504.045 1.525 ;
        RECT 503.715 -0.165 504.045 0.165 ;
        RECT 503.72 -0.165 504.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 505.075 1.195 505.405 1.525 ;
        RECT 505.075 -0.165 505.405 0.165 ;
        RECT 505.08 -0.165 505.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 506.435 1.195 506.765 1.525 ;
        RECT 506.435 -0.165 506.765 0.165 ;
        RECT 506.44 -0.165 506.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 507.795 1.195 508.125 1.525 ;
        RECT 507.795 -0.165 508.125 0.165 ;
        RECT 507.8 -0.165 508.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 509.155 1.195 509.485 1.525 ;
        RECT 509.155 -0.165 509.485 0.165 ;
        RECT 509.16 -0.165 509.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 510.515 1.195 510.845 1.525 ;
        RECT 510.515 -0.165 510.845 0.165 ;
        RECT 510.52 -0.165 510.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 511.875 1.195 512.205 1.525 ;
        RECT 511.875 -0.165 512.205 0.165 ;
        RECT 511.88 -0.165 512.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 513.235 1.195 513.565 1.525 ;
        RECT 513.235 -0.165 513.565 0.165 ;
        RECT 513.24 -0.165 513.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 514.595 1.195 514.925 1.525 ;
        RECT 514.595 -0.165 514.925 0.165 ;
        RECT 514.6 -0.165 514.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 515.955 1.195 516.285 1.525 ;
        RECT 515.955 -0.165 516.285 0.165 ;
        RECT 515.96 -0.165 516.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 517.315 1.195 517.645 1.525 ;
        RECT 517.315 -0.165 517.645 0.165 ;
        RECT 517.32 -0.165 517.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 518.675 1.195 519.005 1.525 ;
        RECT 518.675 -0.165 519.005 0.165 ;
        RECT 518.68 -0.165 519 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 520.035 1.195 520.365 1.525 ;
        RECT 520.035 -0.165 520.365 0.165 ;
        RECT 520.04 -0.165 520.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 521.395 1.195 521.725 1.525 ;
        RECT 521.395 -0.165 521.725 0.165 ;
        RECT 521.4 -0.165 521.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 522.755 1.195 523.085 1.525 ;
        RECT 522.755 -0.165 523.085 0.165 ;
        RECT 522.76 -0.165 523.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 524.115 1.195 524.445 1.525 ;
        RECT 524.115 -0.165 524.445 0.165 ;
        RECT 524.12 -0.165 524.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 525.475 1.195 525.805 1.525 ;
        RECT 525.475 -0.165 525.805 0.165 ;
        RECT 525.48 -0.165 525.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 526.835 1.195 527.165 1.525 ;
        RECT 526.835 -0.165 527.165 0.165 ;
        RECT 526.84 -0.165 527.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 528.195 1.195 528.525 1.525 ;
        RECT 528.195 -0.165 528.525 0.165 ;
        RECT 528.2 -0.165 528.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 529.555 1.195 529.885 1.525 ;
        RECT 529.555 -0.165 529.885 0.165 ;
        RECT 529.56 -0.165 529.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 530.915 1.195 531.245 1.525 ;
        RECT 530.915 -0.165 531.245 0.165 ;
        RECT 530.92 -0.165 531.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 532.275 1.195 532.605 1.525 ;
        RECT 532.275 -0.165 532.605 0.165 ;
        RECT 532.28 -0.165 532.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 533.635 1.195 533.965 1.525 ;
        RECT 533.635 -0.165 533.965 0.165 ;
        RECT 533.64 -0.165 533.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 534.995 1.195 535.325 1.525 ;
        RECT 534.995 -0.165 535.325 0.165 ;
        RECT 535 -0.165 535.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 536.355 1.195 536.685 1.525 ;
        RECT 536.355 -0.165 536.685 0.165 ;
        RECT 536.36 -0.165 536.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 537.715 1.195 538.045 1.525 ;
        RECT 537.715 -0.165 538.045 0.165 ;
        RECT 537.72 -0.165 538.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 539.075 1.195 539.405 1.525 ;
        RECT 539.075 -0.165 539.405 0.165 ;
        RECT 539.08 -0.165 539.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 540.435 1.195 540.765 1.525 ;
        RECT 540.435 -0.165 540.765 0.165 ;
        RECT 540.44 -0.165 540.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 541.795 1.195 542.125 1.525 ;
        RECT 541.795 -0.165 542.125 0.165 ;
        RECT 541.8 -0.165 542.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 543.155 1.195 543.485 1.525 ;
        RECT 543.155 -0.165 543.485 0.165 ;
        RECT 543.16 -0.165 543.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 544.515 1.195 544.845 1.525 ;
        RECT 544.515 -0.165 544.845 0.165 ;
        RECT 544.52 -0.165 544.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 545.875 1.195 546.205 1.525 ;
        RECT 545.875 -0.165 546.205 0.165 ;
        RECT 545.88 -0.165 546.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 547.235 1.195 547.565 1.525 ;
        RECT 547.235 -0.165 547.565 0.165 ;
        RECT 547.24 -0.165 547.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 548.595 1.195 548.925 1.525 ;
        RECT 548.595 -0.165 548.925 0.165 ;
        RECT 548.6 -0.165 548.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 549.955 1.195 550.285 1.525 ;
        RECT 549.955 -0.165 550.285 0.165 ;
        RECT 549.96 -0.165 550.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 551.315 1.195 551.645 1.525 ;
        RECT 551.315 -0.165 551.645 0.165 ;
        RECT 551.32 -0.165 551.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 552.675 1.195 553.005 1.525 ;
        RECT 552.675 -0.165 553.005 0.165 ;
        RECT 552.68 -0.165 553 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 554.035 1.195 554.365 1.525 ;
        RECT 554.035 -0.165 554.365 0.165 ;
        RECT 554.04 -0.165 554.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 555.395 1.195 555.725 1.525 ;
        RECT 555.395 -0.165 555.725 0.165 ;
        RECT 555.4 -0.165 555.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 556.755 1.195 557.085 1.525 ;
        RECT 556.755 -0.165 557.085 0.165 ;
        RECT 556.76 -0.165 557.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 558.115 1.195 558.445 1.525 ;
        RECT 558.115 -0.165 558.445 0.165 ;
        RECT 558.12 -0.165 558.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 559.475 1.195 559.805 1.525 ;
        RECT 559.475 -0.165 559.805 0.165 ;
        RECT 559.48 -0.165 559.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 560.835 1.195 561.165 1.525 ;
        RECT 560.835 -0.165 561.165 0.165 ;
        RECT 560.84 -0.165 561.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 562.195 1.195 562.525 1.525 ;
        RECT 562.195 -0.165 562.525 0.165 ;
        RECT 562.2 -0.165 562.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 563.555 1.195 563.885 1.525 ;
        RECT 563.555 -0.165 563.885 0.165 ;
        RECT 563.56 -0.165 563.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 564.915 1.195 565.245 1.525 ;
        RECT 564.915 -0.165 565.245 0.165 ;
        RECT 564.92 -0.165 565.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 566.275 1.195 566.605 1.525 ;
        RECT 566.275 -0.165 566.605 0.165 ;
        RECT 566.28 -0.165 566.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 567.635 1.195 567.965 1.525 ;
        RECT 567.635 -0.165 567.965 0.165 ;
        RECT 567.64 -0.165 567.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 568.995 1.195 569.325 1.525 ;
        RECT 568.995 -0.165 569.325 0.165 ;
        RECT 569 -0.165 569.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 570.355 1.195 570.685 1.525 ;
        RECT 570.355 -0.165 570.685 0.165 ;
        RECT 570.36 -0.165 570.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 571.715 1.195 572.045 1.525 ;
        RECT 571.715 -0.165 572.045 0.165 ;
        RECT 571.72 -0.165 572.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 573.075 1.195 573.405 1.525 ;
        RECT 573.075 -0.165 573.405 0.165 ;
        RECT 573.08 -0.165 573.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 574.435 1.195 574.765 1.525 ;
        RECT 574.435 -0.165 574.765 0.165 ;
        RECT 574.44 -0.165 574.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 575.795 1.195 576.125 1.525 ;
        RECT 575.795 -0.165 576.125 0.165 ;
        RECT 575.8 -0.165 576.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 577.155 1.195 577.485 1.525 ;
        RECT 577.155 -0.165 577.485 0.165 ;
        RECT 577.16 -0.165 577.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 578.515 1.195 578.845 1.525 ;
        RECT 578.515 -0.165 578.845 0.165 ;
        RECT 578.52 -0.165 578.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 579.875 1.195 580.205 1.525 ;
        RECT 579.875 -0.165 580.205 0.165 ;
        RECT 579.88 -0.165 580.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 581.235 1.195 581.565 1.525 ;
        RECT 581.235 -0.165 581.565 0.165 ;
        RECT 581.24 -0.165 581.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 582.595 1.195 582.925 1.525 ;
        RECT 582.595 -0.165 582.925 0.165 ;
        RECT 582.6 -0.165 582.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 583.955 1.195 584.285 1.525 ;
        RECT 583.955 -0.165 584.285 0.165 ;
        RECT 583.96 -0.165 584.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 585.315 1.195 585.645 1.525 ;
        RECT 585.315 -0.165 585.645 0.165 ;
        RECT 585.32 -0.165 585.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 586.675 1.195 587.005 1.525 ;
        RECT 586.675 -0.165 587.005 0.165 ;
        RECT 586.68 -0.165 587 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 588.035 1.195 588.365 1.525 ;
        RECT 588.035 -0.165 588.365 0.165 ;
        RECT 588.04 -0.165 588.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 589.395 1.195 589.725 1.525 ;
        RECT 589.395 -0.165 589.725 0.165 ;
        RECT 589.4 -0.165 589.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 590.755 1.195 591.085 1.525 ;
        RECT 590.755 -0.165 591.085 0.165 ;
        RECT 590.76 -0.165 591.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 592.115 1.195 592.445 1.525 ;
        RECT 592.115 -0.165 592.445 0.165 ;
        RECT 592.12 -0.165 592.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 593.475 1.195 593.805 1.525 ;
        RECT 593.475 -0.165 593.805 0.165 ;
        RECT 593.48 -0.165 593.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 594.835 1.195 595.165 1.525 ;
        RECT 594.835 -0.165 595.165 0.165 ;
        RECT 594.84 -0.165 595.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 596.195 1.195 596.525 1.525 ;
        RECT 596.195 -0.165 596.525 0.165 ;
        RECT 596.2 -0.165 596.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 597.555 1.195 597.885 1.525 ;
        RECT 597.555 -0.165 597.885 0.165 ;
        RECT 597.56 -0.165 597.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 598.915 1.195 599.245 1.525 ;
        RECT 598.915 -0.165 599.245 0.165 ;
        RECT 598.92 -0.165 599.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 600.275 1.195 600.605 1.525 ;
        RECT 600.275 -0.165 600.605 0.165 ;
        RECT 600.28 -0.165 600.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 601.635 1.195 601.965 1.525 ;
        RECT 601.635 -0.165 601.965 0.165 ;
        RECT 601.64 -0.165 601.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 602.995 1.195 603.325 1.525 ;
        RECT 602.995 -0.165 603.325 0.165 ;
        RECT 603 -0.165 603.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 604.355 1.195 604.685 1.525 ;
        RECT 604.355 -0.165 604.685 0.165 ;
        RECT 604.36 -0.165 604.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 605.715 1.195 606.045 1.525 ;
        RECT 605.715 -0.165 606.045 0.165 ;
        RECT 605.72 -0.165 606.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 607.075 1.195 607.405 1.525 ;
        RECT 607.075 -0.165 607.405 0.165 ;
        RECT 607.08 -0.165 607.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 608.435 1.195 608.765 1.525 ;
        RECT 608.435 -0.165 608.765 0.165 ;
        RECT 608.44 -0.165 608.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 609.795 1.195 610.125 1.525 ;
        RECT 609.795 -0.165 610.125 0.165 ;
        RECT 609.8 -0.165 610.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 611.155 1.195 611.485 1.525 ;
        RECT 611.155 -0.165 611.485 0.165 ;
        RECT 611.16 -0.165 611.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 612.515 1.195 612.845 1.525 ;
        RECT 612.515 -0.165 612.845 0.165 ;
        RECT 612.52 -0.165 612.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 613.875 1.195 614.205 1.525 ;
        RECT 613.875 -0.165 614.205 0.165 ;
        RECT 613.88 -0.165 614.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 615.235 1.195 615.565 1.525 ;
        RECT 615.235 -0.165 615.565 0.165 ;
        RECT 615.24 -0.165 615.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 616.595 1.195 616.925 1.525 ;
        RECT 616.595 -0.165 616.925 0.165 ;
        RECT 616.6 -0.165 616.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 617.955 1.195 618.285 1.525 ;
        RECT 617.955 -0.165 618.285 0.165 ;
        RECT 617.96 -0.165 618.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 619.315 1.195 619.645 1.525 ;
        RECT 619.315 -0.165 619.645 0.165 ;
        RECT 619.32 -0.165 619.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 620.675 1.195 621.005 1.525 ;
        RECT 620.675 -0.165 621.005 0.165 ;
        RECT 620.68 -0.165 621 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 622.035 1.195 622.365 1.525 ;
        RECT 622.035 -0.165 622.365 0.165 ;
        RECT 622.04 -0.165 622.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 623.395 1.195 623.725 1.525 ;
        RECT 623.395 -0.165 623.725 0.165 ;
        RECT 623.4 -0.165 623.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 624.755 1.195 625.085 1.525 ;
        RECT 624.755 -0.165 625.085 0.165 ;
        RECT 624.76 -0.165 625.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 626.115 1.195 626.445 1.525 ;
        RECT 626.115 -0.165 626.445 0.165 ;
        RECT 626.12 -0.165 626.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 627.475 1.195 627.805 1.525 ;
        RECT 627.475 -0.165 627.805 0.165 ;
        RECT 627.48 -0.165 627.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 628.835 1.195 629.165 1.525 ;
        RECT 628.835 -0.165 629.165 0.165 ;
        RECT 628.84 -0.165 629.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 630.195 1.195 630.525 1.525 ;
        RECT 630.195 -0.165 630.525 0.165 ;
        RECT 630.2 -0.165 630.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 631.555 1.195 631.885 1.525 ;
        RECT 631.555 -0.165 631.885 0.165 ;
        RECT 631.56 -0.165 631.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 632.915 1.195 633.245 1.525 ;
        RECT 632.915 -0.165 633.245 0.165 ;
        RECT 632.92 -0.165 633.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 634.275 1.195 634.605 1.525 ;
        RECT 634.275 -0.165 634.605 0.165 ;
        RECT 634.28 -0.165 634.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 635.635 1.195 635.965 1.525 ;
        RECT 635.635 -0.165 635.965 0.165 ;
        RECT 635.64 -0.165 635.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 636.995 1.195 637.325 1.525 ;
        RECT 636.995 -0.165 637.325 0.165 ;
        RECT 637 -0.165 637.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 638.355 1.195 638.685 1.525 ;
        RECT 638.355 -0.165 638.685 0.165 ;
        RECT 638.36 -0.165 638.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 639.715 1.195 640.045 1.525 ;
        RECT 639.715 -0.165 640.045 0.165 ;
        RECT 639.72 -0.165 640.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 641.075 1.195 641.405 1.525 ;
        RECT 641.075 -0.165 641.405 0.165 ;
        RECT 641.08 -0.165 641.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 642.435 1.195 642.765 1.525 ;
        RECT 642.435 -0.165 642.765 0.165 ;
        RECT 642.44 -0.165 642.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 643.795 1.195 644.125 1.525 ;
        RECT 643.795 -0.165 644.125 0.165 ;
        RECT 643.8 -0.165 644.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 645.155 1.195 645.485 1.525 ;
        RECT 645.155 -0.165 645.485 0.165 ;
        RECT 645.16 -0.165 645.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 646.515 1.195 646.845 1.525 ;
        RECT 646.515 -0.165 646.845 0.165 ;
        RECT 646.52 -0.165 646.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 647.875 1.195 648.205 1.525 ;
        RECT 647.875 -0.165 648.205 0.165 ;
        RECT 647.88 -0.165 648.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 649.235 1.195 649.565 1.525 ;
        RECT 649.235 -0.165 649.565 0.165 ;
        RECT 649.24 -0.165 649.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 650.595 1.195 650.925 1.525 ;
        RECT 650.595 -0.165 650.925 0.165 ;
        RECT 650.6 -0.165 650.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 651.955 1.195 652.285 1.525 ;
        RECT 651.955 -0.165 652.285 0.165 ;
        RECT 651.96 -0.165 652.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 653.315 1.195 653.645 1.525 ;
        RECT 653.315 -0.165 653.645 0.165 ;
        RECT 653.32 -0.165 653.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 654.675 1.195 655.005 1.525 ;
        RECT 654.675 -0.165 655.005 0.165 ;
        RECT 654.68 -0.165 655 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 656.035 1.195 656.365 1.525 ;
        RECT 656.035 -0.165 656.365 0.165 ;
        RECT 656.04 -0.165 656.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 657.395 1.195 657.725 1.525 ;
        RECT 657.395 -0.165 657.725 0.165 ;
        RECT 657.4 -0.165 657.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 658.755 1.195 659.085 1.525 ;
        RECT 658.755 -0.165 659.085 0.165 ;
        RECT 658.76 -0.165 659.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 660.115 1.195 660.445 1.525 ;
        RECT 660.115 -0.165 660.445 0.165 ;
        RECT 660.12 -0.165 660.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 661.475 1.195 661.805 1.525 ;
        RECT 661.475 -0.165 661.805 0.165 ;
        RECT 661.48 -0.165 661.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 662.835 1.195 663.165 1.525 ;
        RECT 662.835 -0.165 663.165 0.165 ;
        RECT 662.84 -0.165 663.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 664.195 1.195 664.525 1.525 ;
        RECT 664.195 -0.165 664.525 0.165 ;
        RECT 664.2 -0.165 664.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 665.555 1.195 665.885 1.525 ;
        RECT 665.555 -0.165 665.885 0.165 ;
        RECT 665.56 -0.165 665.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 666.915 1.195 667.245 1.525 ;
        RECT 666.915 -0.165 667.245 0.165 ;
        RECT 666.92 -0.165 667.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 668.275 1.195 668.605 1.525 ;
        RECT 668.275 -0.165 668.605 0.165 ;
        RECT 668.28 -0.165 668.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 669.635 1.195 669.965 1.525 ;
        RECT 669.635 -0.165 669.965 0.165 ;
        RECT 669.64 -0.165 669.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 670.995 1.195 671.325 1.525 ;
        RECT 670.995 -0.165 671.325 0.165 ;
        RECT 671 -0.165 671.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 672.355 1.195 672.685 1.525 ;
        RECT 672.355 -0.165 672.685 0.165 ;
        RECT 672.36 -0.165 672.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 673.715 1.195 674.045 1.525 ;
        RECT 673.715 -0.165 674.045 0.165 ;
        RECT 673.72 -0.165 674.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 675.075 1.195 675.405 1.525 ;
        RECT 675.075 -0.165 675.405 0.165 ;
        RECT 675.08 -0.165 675.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 676.435 1.195 676.765 1.525 ;
        RECT 676.435 -0.165 676.765 0.165 ;
        RECT 676.44 -0.165 676.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 677.795 1.195 678.125 1.525 ;
        RECT 677.795 -0.165 678.125 0.165 ;
        RECT 677.8 -0.165 678.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 679.155 1.195 679.485 1.525 ;
        RECT 679.155 -0.165 679.485 0.165 ;
        RECT 679.16 -0.165 679.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 680.515 1.195 680.845 1.525 ;
        RECT 680.515 -0.165 680.845 0.165 ;
        RECT 680.52 -0.165 680.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 681.875 1.195 682.205 1.525 ;
        RECT 681.875 -0.165 682.205 0.165 ;
        RECT 681.88 -0.165 682.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 683.235 1.195 683.565 1.525 ;
        RECT 683.235 -0.165 683.565 0.165 ;
        RECT 683.24 -0.165 683.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 684.595 1.195 684.925 1.525 ;
        RECT 684.595 -0.165 684.925 0.165 ;
        RECT 684.6 -0.165 684.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 685.955 1.195 686.285 1.525 ;
        RECT 685.955 -0.165 686.285 0.165 ;
        RECT 685.96 -0.165 686.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 687.315 1.195 687.645 1.525 ;
        RECT 687.315 -0.165 687.645 0.165 ;
        RECT 687.32 -0.165 687.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 688.675 1.195 689.005 1.525 ;
        RECT 688.675 -0.165 689.005 0.165 ;
        RECT 688.68 -0.165 689 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 690.035 1.195 690.365 1.525 ;
        RECT 690.035 -0.165 690.365 0.165 ;
        RECT 690.04 -0.165 690.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 691.395 1.195 691.725 1.525 ;
        RECT 691.395 -0.165 691.725 0.165 ;
        RECT 691.4 -0.165 691.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 692.755 1.195 693.085 1.525 ;
        RECT 692.755 -0.165 693.085 0.165 ;
        RECT 692.76 -0.165 693.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 694.115 1.195 694.445 1.525 ;
        RECT 694.115 -0.165 694.445 0.165 ;
        RECT 694.12 -0.165 694.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 695.475 1.195 695.805 1.525 ;
        RECT 695.475 -0.165 695.805 0.165 ;
        RECT 695.48 -0.165 695.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 696.835 1.195 697.165 1.525 ;
        RECT 696.835 -0.165 697.165 0.165 ;
        RECT 696.84 -0.165 697.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 698.195 1.195 698.525 1.525 ;
        RECT 698.195 -0.165 698.525 0.165 ;
        RECT 698.2 -0.165 698.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 699.555 1.195 699.885 1.525 ;
        RECT 699.555 -0.165 699.885 0.165 ;
        RECT 699.56 -0.165 699.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 700.915 1.195 701.245 1.525 ;
        RECT 700.915 -0.165 701.245 0.165 ;
        RECT 700.92 -0.165 701.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 702.275 1.195 702.605 1.525 ;
        RECT 702.275 -0.165 702.605 0.165 ;
        RECT 702.28 -0.165 702.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 703.635 1.195 703.965 1.525 ;
        RECT 703.635 -0.165 703.965 0.165 ;
        RECT 703.64 -0.165 703.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 704.995 1.195 705.325 1.525 ;
        RECT 704.995 -0.165 705.325 0.165 ;
        RECT 705 -0.165 705.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 706.355 1.195 706.685 1.525 ;
        RECT 706.355 -0.165 706.685 0.165 ;
        RECT 706.36 -0.165 706.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 707.715 1.195 708.045 1.525 ;
        RECT 707.715 -0.165 708.045 0.165 ;
        RECT 707.72 -0.165 708.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 709.075 1.195 709.405 1.525 ;
        RECT 709.075 -0.165 709.405 0.165 ;
        RECT 709.08 -0.165 709.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 710.435 1.195 710.765 1.525 ;
        RECT 710.435 -0.165 710.765 0.165 ;
        RECT 710.44 -0.165 710.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 711.795 1.195 712.125 1.525 ;
        RECT 711.795 -0.165 712.125 0.165 ;
        RECT 711.8 -0.165 712.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 713.155 1.195 713.485 1.525 ;
        RECT 713.155 -0.165 713.485 0.165 ;
        RECT 713.16 -0.165 713.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 714.515 1.195 714.845 1.525 ;
        RECT 714.515 -0.165 714.845 0.165 ;
        RECT 714.52 -0.165 714.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 715.875 1.195 716.205 1.525 ;
        RECT 715.875 -0.165 716.205 0.165 ;
        RECT 715.88 -0.165 716.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 717.235 1.195 717.565 1.525 ;
        RECT 717.235 -0.165 717.565 0.165 ;
        RECT 717.24 -0.165 717.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 718.595 1.195 718.925 1.525 ;
        RECT 718.595 -0.165 718.925 0.165 ;
        RECT 718.6 -0.165 718.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 719.955 1.195 720.285 1.525 ;
        RECT 719.955 -0.165 720.285 0.165 ;
        RECT 719.96 -0.165 720.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 721.315 1.195 721.645 1.525 ;
        RECT 721.315 -0.165 721.645 0.165 ;
        RECT 721.32 -0.165 721.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 722.675 1.195 723.005 1.525 ;
        RECT 722.675 -0.165 723.005 0.165 ;
        RECT 722.68 -0.165 723 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 724.035 1.195 724.365 1.525 ;
        RECT 724.035 -0.165 724.365 0.165 ;
        RECT 724.04 -0.165 724.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 725.395 1.195 725.725 1.525 ;
        RECT 725.395 -0.165 725.725 0.165 ;
        RECT 725.4 -0.165 725.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 726.755 1.195 727.085 1.525 ;
        RECT 726.755 -0.165 727.085 0.165 ;
        RECT 726.76 -0.165 727.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 728.115 1.195 728.445 1.525 ;
        RECT 728.115 -0.165 728.445 0.165 ;
        RECT 728.12 -0.165 728.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 729.475 1.195 729.805 1.525 ;
        RECT 729.475 -0.165 729.805 0.165 ;
        RECT 729.48 -0.165 729.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 730.835 1.195 731.165 1.525 ;
        RECT 730.835 -0.165 731.165 0.165 ;
        RECT 730.84 -0.165 731.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 732.195 1.195 732.525 1.525 ;
        RECT 732.195 -0.165 732.525 0.165 ;
        RECT 732.2 -0.165 732.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 733.555 1.195 733.885 1.525 ;
        RECT 733.555 -0.165 733.885 0.165 ;
        RECT 733.56 -0.165 733.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 734.915 1.195 735.245 1.525 ;
        RECT 734.915 -0.165 735.245 0.165 ;
        RECT 734.92 -0.165 735.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 736.275 1.195 736.605 1.525 ;
        RECT 736.275 -0.165 736.605 0.165 ;
        RECT 736.28 -0.165 736.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 737.635 1.195 737.965 1.525 ;
        RECT 737.635 -0.165 737.965 0.165 ;
        RECT 737.64 -0.165 737.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 738.995 1.195 739.325 1.525 ;
        RECT 738.995 -0.165 739.325 0.165 ;
        RECT 739 -0.165 739.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 740.355 1.195 740.685 1.525 ;
        RECT 740.355 -0.165 740.685 0.165 ;
        RECT 740.36 -0.165 740.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 741.715 1.195 742.045 1.525 ;
        RECT 741.715 -0.165 742.045 0.165 ;
        RECT 741.72 -0.165 742.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 743.075 1.195 743.405 1.525 ;
        RECT 743.075 -0.165 743.405 0.165 ;
        RECT 743.08 -0.165 743.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 744.435 1.195 744.765 1.525 ;
        RECT 744.435 -0.165 744.765 0.165 ;
        RECT 744.44 -0.165 744.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 745.795 1.195 746.125 1.525 ;
        RECT 745.795 -0.165 746.125 0.165 ;
        RECT 745.8 -0.165 746.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 747.155 1.195 747.485 1.525 ;
        RECT 747.155 -0.165 747.485 0.165 ;
        RECT 747.16 -0.165 747.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 748.515 1.195 748.845 1.525 ;
        RECT 748.515 -0.165 748.845 0.165 ;
        RECT 748.52 -0.165 748.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 749.875 1.195 750.205 1.525 ;
        RECT 749.875 -0.165 750.205 0.165 ;
        RECT 749.88 -0.165 750.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 751.235 1.195 751.565 1.525 ;
        RECT 751.235 -0.165 751.565 0.165 ;
        RECT 751.24 -0.165 751.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 752.595 1.195 752.925 1.525 ;
        RECT 752.595 -0.165 752.925 0.165 ;
        RECT 752.6 -0.165 752.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 753.955 1.195 754.285 1.525 ;
        RECT 753.955 -0.165 754.285 0.165 ;
        RECT 753.96 -0.165 754.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 755.315 1.195 755.645 1.525 ;
        RECT 755.315 -0.165 755.645 0.165 ;
        RECT 755.32 -0.165 755.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 756.675 1.195 757.005 1.525 ;
        RECT 756.675 -0.165 757.005 0.165 ;
        RECT 756.68 -0.165 757 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 758.035 1.195 758.365 1.525 ;
        RECT 758.035 -0.165 758.365 0.165 ;
        RECT 758.04 -0.165 758.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 759.395 1.195 759.725 1.525 ;
        RECT 759.395 -0.165 759.725 0.165 ;
        RECT 759.4 -0.165 759.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 760.755 1.195 761.085 1.525 ;
        RECT 760.755 -0.165 761.085 0.165 ;
        RECT 760.76 -0.165 761.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 762.115 1.195 762.445 1.525 ;
        RECT 762.115 -0.165 762.445 0.165 ;
        RECT 762.12 -0.165 762.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 763.475 3.915 763.805 4.245 ;
        RECT 763.475 1.195 763.805 1.525 ;
        RECT 763.475 -0.165 763.805 0.165 ;
        RECT 763.48 -0.165 763.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 764.835 3.915 765.165 4.245 ;
        RECT 764.835 1.195 765.165 1.525 ;
        RECT 764.835 -0.165 765.165 0.165 ;
        RECT 764.84 -0.165 765.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 766.195 3.915 766.525 4.245 ;
        RECT 766.195 2.555 766.525 2.885 ;
        RECT 766.195 1.195 766.525 1.525 ;
        RECT 766.195 -0.165 766.525 0.165 ;
        RECT 766.2 -0.165 766.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 767.555 3.915 767.885 4.245 ;
        RECT 767.555 2.555 767.885 2.885 ;
        RECT 767.555 1.195 767.885 1.525 ;
        RECT 767.555 -0.165 767.885 0.165 ;
        RECT 767.56 -0.165 767.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 768.915 5.275 769.245 5.605 ;
        RECT 768.915 3.915 769.245 4.245 ;
        RECT 768.915 2.555 769.245 2.885 ;
        RECT 768.915 1.195 769.245 1.525 ;
        RECT 768.915 -0.165 769.245 0.165 ;
        RECT 768.92 -0.165 769.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -2.205 5.275 -1.875 5.605 ;
        RECT -2.205 3.915 -1.875 4.245 ;
        RECT -2.205 2.555 -1.875 2.885 ;
        RECT -2.205 1.195 -1.875 1.525 ;
        RECT -2.205 -0.165 -1.875 0.165 ;
        RECT -2.2 -0.165 -1.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.845 5.275 -0.515 5.605 ;
        RECT -0.845 3.915 -0.515 4.245 ;
        RECT -0.845 2.555 -0.515 2.885 ;
        RECT -0.845 1.195 -0.515 1.525 ;
        RECT -0.845 -0.165 -0.515 0.165 ;
        RECT -0.84 -0.165 -0.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.515 3.915 0.845 4.245 ;
        RECT 0.515 2.555 0.845 2.885 ;
        RECT 0.515 1.195 0.845 1.525 ;
        RECT 0.515 -0.165 0.845 0.165 ;
        RECT 0.52 -0.165 0.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.875 3.915 2.205 4.245 ;
        RECT 1.875 1.195 2.205 1.525 ;
        RECT 1.875 -0.165 2.205 0.165 ;
        RECT 1.88 -0.165 2.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.235 3.915 3.565 4.245 ;
        RECT 3.235 1.195 3.565 1.525 ;
        RECT 3.235 -0.165 3.565 0.165 ;
        RECT 3.24 -0.165 3.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.595 1.195 4.925 1.525 ;
        RECT 4.595 -0.165 4.925 0.165 ;
        RECT 4.6 -0.165 4.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.955 1.195 6.285 1.525 ;
        RECT 5.955 -0.165 6.285 0.165 ;
        RECT 5.96 -0.165 6.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.315 1.195 7.645 1.525 ;
        RECT 7.315 -0.165 7.645 0.165 ;
        RECT 7.32 -0.165 7.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.675 1.195 9.005 1.525 ;
        RECT 8.675 -0.165 9.005 0.165 ;
        RECT 8.68 -0.165 9 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.035 1.195 10.365 1.525 ;
        RECT 10.035 -0.165 10.365 0.165 ;
        RECT 10.04 -0.165 10.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.395 1.195 11.725 1.525 ;
        RECT 11.395 -0.165 11.725 0.165 ;
        RECT 11.4 -0.165 11.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.755 1.195 13.085 1.525 ;
        RECT 12.755 -0.165 13.085 0.165 ;
        RECT 12.76 -0.165 13.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.115 1.195 14.445 1.525 ;
        RECT 14.115 -0.165 14.445 0.165 ;
        RECT 14.12 -0.165 14.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.475 1.195 15.805 1.525 ;
        RECT 15.475 -0.165 15.805 0.165 ;
        RECT 15.48 -0.165 15.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.835 1.195 17.165 1.525 ;
        RECT 16.835 -0.165 17.165 0.165 ;
        RECT 16.84 -0.165 17.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.195 1.195 18.525 1.525 ;
        RECT 18.195 -0.165 18.525 0.165 ;
        RECT 18.2 -0.165 18.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.555 1.195 19.885 1.525 ;
        RECT 19.555 -0.165 19.885 0.165 ;
        RECT 19.56 -0.165 19.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.915 1.195 21.245 1.525 ;
        RECT 20.915 -0.165 21.245 0.165 ;
        RECT 20.92 -0.165 21.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.275 1.195 22.605 1.525 ;
        RECT 22.275 -0.165 22.605 0.165 ;
        RECT 22.28 -0.165 22.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.635 1.195 23.965 1.525 ;
        RECT 23.635 -0.165 23.965 0.165 ;
        RECT 23.64 -0.165 23.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.995 1.195 25.325 1.525 ;
        RECT 24.995 -0.165 25.325 0.165 ;
        RECT 25 -0.165 25.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.355 1.195 26.685 1.525 ;
        RECT 26.355 -0.165 26.685 0.165 ;
        RECT 26.36 -0.165 26.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.715 1.195 28.045 1.525 ;
        RECT 27.715 -0.165 28.045 0.165 ;
        RECT 27.72 -0.165 28.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.075 1.195 29.405 1.525 ;
        RECT 29.075 -0.165 29.405 0.165 ;
        RECT 29.08 -0.165 29.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.435 1.195 30.765 1.525 ;
        RECT 30.435 -0.165 30.765 0.165 ;
        RECT 30.44 -0.165 30.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.795 1.195 32.125 1.525 ;
        RECT 31.795 -0.165 32.125 0.165 ;
        RECT 31.8 -0.165 32.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.155 1.195 33.485 1.525 ;
        RECT 33.155 -0.165 33.485 0.165 ;
        RECT 33.16 -0.165 33.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.515 1.195 34.845 1.525 ;
        RECT 34.515 -0.165 34.845 0.165 ;
        RECT 34.52 -0.165 34.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.875 1.195 36.205 1.525 ;
        RECT 35.875 -0.165 36.205 0.165 ;
        RECT 35.88 -0.165 36.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.235 1.195 37.565 1.525 ;
        RECT 37.235 -0.165 37.565 0.165 ;
        RECT 37.24 -0.165 37.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.595 1.195 38.925 1.525 ;
        RECT 38.595 -0.165 38.925 0.165 ;
        RECT 38.6 -0.165 38.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.955 1.195 40.285 1.525 ;
        RECT 39.955 -0.165 40.285 0.165 ;
        RECT 39.96 -0.165 40.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.315 1.195 41.645 1.525 ;
        RECT 41.315 -0.165 41.645 0.165 ;
        RECT 41.32 -0.165 41.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.675 1.195 43.005 1.525 ;
        RECT 42.675 -0.165 43.005 0.165 ;
        RECT 42.68 -0.165 43 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.035 1.195 44.365 1.525 ;
        RECT 44.035 -0.165 44.365 0.165 ;
        RECT 44.04 -0.165 44.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.395 1.195 45.725 1.525 ;
        RECT 45.395 -0.165 45.725 0.165 ;
        RECT 45.4 -0.165 45.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.755 1.195 47.085 1.525 ;
        RECT 46.755 -0.165 47.085 0.165 ;
        RECT 46.76 -0.165 47.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.115 1.195 48.445 1.525 ;
        RECT 48.115 -0.165 48.445 0.165 ;
        RECT 48.12 -0.165 48.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.475 1.195 49.805 1.525 ;
        RECT 49.475 -0.165 49.805 0.165 ;
        RECT 49.48 -0.165 49.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.835 1.195 51.165 1.525 ;
        RECT 50.835 -0.165 51.165 0.165 ;
        RECT 50.84 -0.165 51.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.195 1.195 52.525 1.525 ;
        RECT 52.195 -0.165 52.525 0.165 ;
        RECT 52.2 -0.165 52.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.555 1.195 53.885 1.525 ;
        RECT 53.555 -0.165 53.885 0.165 ;
        RECT 53.56 -0.165 53.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.915 1.195 55.245 1.525 ;
        RECT 54.915 -0.165 55.245 0.165 ;
        RECT 54.92 -0.165 55.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.275 1.195 56.605 1.525 ;
        RECT 56.275 -0.165 56.605 0.165 ;
        RECT 56.28 -0.165 56.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.635 1.195 57.965 1.525 ;
        RECT 57.635 -0.165 57.965 0.165 ;
        RECT 57.64 -0.165 57.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.995 1.195 59.325 1.525 ;
        RECT 58.995 -0.165 59.325 0.165 ;
        RECT 59 -0.165 59.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.355 1.195 60.685 1.525 ;
        RECT 60.355 -0.165 60.685 0.165 ;
        RECT 60.36 -0.165 60.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.715 1.195 62.045 1.525 ;
        RECT 61.715 -0.165 62.045 0.165 ;
        RECT 61.72 -0.165 62.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.075 1.195 63.405 1.525 ;
        RECT 63.075 -0.165 63.405 0.165 ;
        RECT 63.08 -0.165 63.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.435 1.195 64.765 1.525 ;
        RECT 64.435 -0.165 64.765 0.165 ;
        RECT 64.44 -0.165 64.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.795 1.195 66.125 1.525 ;
        RECT 65.795 -0.165 66.125 0.165 ;
        RECT 65.8 -0.165 66.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.155 1.195 67.485 1.525 ;
        RECT 67.155 -0.165 67.485 0.165 ;
        RECT 67.16 -0.165 67.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.515 1.195 68.845 1.525 ;
        RECT 68.515 -0.165 68.845 0.165 ;
        RECT 68.52 -0.165 68.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.875 1.195 70.205 1.525 ;
        RECT 69.875 -0.165 70.205 0.165 ;
        RECT 69.88 -0.165 70.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.235 1.195 71.565 1.525 ;
        RECT 71.235 -0.165 71.565 0.165 ;
        RECT 71.24 -0.165 71.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.595 1.195 72.925 1.525 ;
        RECT 72.595 -0.165 72.925 0.165 ;
        RECT 72.6 -0.165 72.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 1.195 74.285 1.525 ;
        RECT 73.955 -0.165 74.285 0.165 ;
        RECT 73.96 -0.165 74.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.315 1.195 75.645 1.525 ;
        RECT 75.315 -0.165 75.645 0.165 ;
        RECT 75.32 -0.165 75.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 76.675 1.195 77.005 1.525 ;
        RECT 76.675 -0.165 77.005 0.165 ;
        RECT 76.68 -0.165 77 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.035 1.195 78.365 1.525 ;
        RECT 78.035 -0.165 78.365 0.165 ;
        RECT 78.04 -0.165 78.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 79.395 1.195 79.725 1.525 ;
        RECT 79.395 -0.165 79.725 0.165 ;
        RECT 79.4 -0.165 79.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.755 1.195 81.085 1.525 ;
        RECT 80.755 -0.165 81.085 0.165 ;
        RECT 80.76 -0.165 81.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.115 1.195 82.445 1.525 ;
        RECT 82.115 -0.165 82.445 0.165 ;
        RECT 82.12 -0.165 82.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 83.475 1.195 83.805 1.525 ;
        RECT 83.475 -0.165 83.805 0.165 ;
        RECT 83.48 -0.165 83.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.835 1.195 85.165 1.525 ;
        RECT 84.835 -0.165 85.165 0.165 ;
        RECT 84.84 -0.165 85.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.195 1.195 86.525 1.525 ;
        RECT 86.195 -0.165 86.525 0.165 ;
        RECT 86.2 -0.165 86.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.555 1.195 87.885 1.525 ;
        RECT 87.555 -0.165 87.885 0.165 ;
        RECT 87.56 -0.165 87.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.915 1.195 89.245 1.525 ;
        RECT 88.915 -0.165 89.245 0.165 ;
        RECT 88.92 -0.165 89.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.275 1.195 90.605 1.525 ;
        RECT 90.275 -0.165 90.605 0.165 ;
        RECT 90.28 -0.165 90.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 91.635 1.195 91.965 1.525 ;
        RECT 91.635 -0.165 91.965 0.165 ;
        RECT 91.64 -0.165 91.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.995 1.195 93.325 1.525 ;
        RECT 92.995 -0.165 93.325 0.165 ;
        RECT 93 -0.165 93.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.355 1.195 94.685 1.525 ;
        RECT 94.355 -0.165 94.685 0.165 ;
        RECT 94.36 -0.165 94.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.715 1.195 96.045 1.525 ;
        RECT 95.715 -0.165 96.045 0.165 ;
        RECT 95.72 -0.165 96.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.075 1.195 97.405 1.525 ;
        RECT 97.075 -0.165 97.405 0.165 ;
        RECT 97.08 -0.165 97.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.435 1.195 98.765 1.525 ;
        RECT 98.435 -0.165 98.765 0.165 ;
        RECT 98.44 -0.165 98.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.795 1.195 100.125 1.525 ;
        RECT 99.795 -0.165 100.125 0.165 ;
        RECT 99.8 -0.165 100.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.155 1.195 101.485 1.525 ;
        RECT 101.155 -0.165 101.485 0.165 ;
        RECT 101.16 -0.165 101.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.515 1.195 102.845 1.525 ;
        RECT 102.515 -0.165 102.845 0.165 ;
        RECT 102.52 -0.165 102.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.875 1.195 104.205 1.525 ;
        RECT 103.875 -0.165 104.205 0.165 ;
        RECT 103.88 -0.165 104.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.235 1.195 105.565 1.525 ;
        RECT 105.235 -0.165 105.565 0.165 ;
        RECT 105.24 -0.165 105.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.595 1.195 106.925 1.525 ;
        RECT 106.595 -0.165 106.925 0.165 ;
        RECT 106.6 -0.165 106.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.955 1.195 108.285 1.525 ;
        RECT 107.955 -0.165 108.285 0.165 ;
        RECT 107.96 -0.165 108.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.315 1.195 109.645 1.525 ;
        RECT 109.315 -0.165 109.645 0.165 ;
        RECT 109.32 -0.165 109.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.675 1.195 111.005 1.525 ;
        RECT 110.675 -0.165 111.005 0.165 ;
        RECT 110.68 -0.165 111 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.035 1.195 112.365 1.525 ;
        RECT 112.035 -0.165 112.365 0.165 ;
        RECT 112.04 -0.165 112.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.395 1.195 113.725 1.525 ;
        RECT 113.395 -0.165 113.725 0.165 ;
        RECT 113.4 -0.165 113.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.755 1.195 115.085 1.525 ;
        RECT 114.755 -0.165 115.085 0.165 ;
        RECT 114.76 -0.165 115.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.115 1.195 116.445 1.525 ;
        RECT 116.115 -0.165 116.445 0.165 ;
        RECT 116.12 -0.165 116.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 117.475 1.195 117.805 1.525 ;
        RECT 117.475 -0.165 117.805 0.165 ;
        RECT 117.48 -0.165 117.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.835 1.195 119.165 1.525 ;
        RECT 118.835 -0.165 119.165 0.165 ;
        RECT 118.84 -0.165 119.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.195 1.195 120.525 1.525 ;
        RECT 120.195 -0.165 120.525 0.165 ;
        RECT 120.2 -0.165 120.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 121.555 1.195 121.885 1.525 ;
        RECT 121.555 -0.165 121.885 0.165 ;
        RECT 121.56 -0.165 121.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.915 1.195 123.245 1.525 ;
        RECT 122.915 -0.165 123.245 0.165 ;
        RECT 122.92 -0.165 123.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.275 1.195 124.605 1.525 ;
        RECT 124.275 -0.165 124.605 0.165 ;
        RECT 124.28 -0.165 124.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.635 1.195 125.965 1.525 ;
        RECT 125.635 -0.165 125.965 0.165 ;
        RECT 125.64 -0.165 125.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.995 1.195 127.325 1.525 ;
        RECT 126.995 -0.165 127.325 0.165 ;
        RECT 127 -0.165 127.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.355 1.195 128.685 1.525 ;
        RECT 128.355 -0.165 128.685 0.165 ;
        RECT 128.36 -0.165 128.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.715 1.195 130.045 1.525 ;
        RECT 129.715 -0.165 130.045 0.165 ;
        RECT 129.72 -0.165 130.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.075 1.195 131.405 1.525 ;
        RECT 131.075 -0.165 131.405 0.165 ;
        RECT 131.08 -0.165 131.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.435 1.195 132.765 1.525 ;
        RECT 132.435 -0.165 132.765 0.165 ;
        RECT 132.44 -0.165 132.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.795 1.195 134.125 1.525 ;
        RECT 133.795 -0.165 134.125 0.165 ;
        RECT 133.8 -0.165 134.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.155 1.195 135.485 1.525 ;
        RECT 135.155 -0.165 135.485 0.165 ;
        RECT 135.16 -0.165 135.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 136.515 1.195 136.845 1.525 ;
        RECT 136.515 -0.165 136.845 0.165 ;
        RECT 136.52 -0.165 136.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.875 1.195 138.205 1.525 ;
        RECT 137.875 -0.165 138.205 0.165 ;
        RECT 137.88 -0.165 138.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.235 1.195 139.565 1.525 ;
        RECT 139.235 -0.165 139.565 0.165 ;
        RECT 139.24 -0.165 139.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.595 1.195 140.925 1.525 ;
        RECT 140.595 -0.165 140.925 0.165 ;
        RECT 140.6 -0.165 140.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.955 1.195 142.285 1.525 ;
        RECT 141.955 -0.165 142.285 0.165 ;
        RECT 141.96 -0.165 142.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.315 1.195 143.645 1.525 ;
        RECT 143.315 -0.165 143.645 0.165 ;
        RECT 143.32 -0.165 143.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 144.675 1.195 145.005 1.525 ;
        RECT 144.675 -0.165 145.005 0.165 ;
        RECT 144.68 -0.165 145 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.035 1.195 146.365 1.525 ;
        RECT 146.035 -0.165 146.365 0.165 ;
        RECT 146.04 -0.165 146.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.395 1.195 147.725 1.525 ;
        RECT 147.395 -0.165 147.725 0.165 ;
        RECT 147.4 -0.165 147.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.755 1.195 149.085 1.525 ;
        RECT 148.755 -0.165 149.085 0.165 ;
        RECT 148.76 -0.165 149.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.115 1.195 150.445 1.525 ;
        RECT 150.115 -0.165 150.445 0.165 ;
        RECT 150.12 -0.165 150.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 151.475 1.195 151.805 1.525 ;
        RECT 151.475 -0.165 151.805 0.165 ;
        RECT 151.48 -0.165 151.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.835 1.195 153.165 1.525 ;
        RECT 152.835 -0.165 153.165 0.165 ;
        RECT 152.84 -0.165 153.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.195 1.195 154.525 1.525 ;
        RECT 154.195 -0.165 154.525 0.165 ;
        RECT 154.2 -0.165 154.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.555 1.195 155.885 1.525 ;
        RECT 155.555 -0.165 155.885 0.165 ;
        RECT 155.56 -0.165 155.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.915 1.195 157.245 1.525 ;
        RECT 156.915 -0.165 157.245 0.165 ;
        RECT 156.92 -0.165 157.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.275 1.195 158.605 1.525 ;
        RECT 158.275 -0.165 158.605 0.165 ;
        RECT 158.28 -0.165 158.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.635 1.195 159.965 1.525 ;
        RECT 159.635 -0.165 159.965 0.165 ;
        RECT 159.64 -0.165 159.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.995 1.195 161.325 1.525 ;
        RECT 160.995 -0.165 161.325 0.165 ;
        RECT 161 -0.165 161.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 162.355 1.195 162.685 1.525 ;
        RECT 162.355 -0.165 162.685 0.165 ;
        RECT 162.36 -0.165 162.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.715 1.195 164.045 1.525 ;
        RECT 163.715 -0.165 164.045 0.165 ;
        RECT 163.72 -0.165 164.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.075 1.195 165.405 1.525 ;
        RECT 165.075 -0.165 165.405 0.165 ;
        RECT 165.08 -0.165 165.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.435 1.195 166.765 1.525 ;
        RECT 166.435 -0.165 166.765 0.165 ;
        RECT 166.44 -0.165 166.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.795 1.195 168.125 1.525 ;
        RECT 167.795 -0.165 168.125 0.165 ;
        RECT 167.8 -0.165 168.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.155 1.195 169.485 1.525 ;
        RECT 169.155 -0.165 169.485 0.165 ;
        RECT 169.16 -0.165 169.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.515 1.195 170.845 1.525 ;
        RECT 170.515 -0.165 170.845 0.165 ;
        RECT 170.52 -0.165 170.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.875 1.195 172.205 1.525 ;
        RECT 171.875 -0.165 172.205 0.165 ;
        RECT 171.88 -0.165 172.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.235 1.195 173.565 1.525 ;
        RECT 173.235 -0.165 173.565 0.165 ;
        RECT 173.24 -0.165 173.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 174.595 1.195 174.925 1.525 ;
        RECT 174.595 -0.165 174.925 0.165 ;
        RECT 174.6 -0.165 174.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.955 1.195 176.285 1.525 ;
        RECT 175.955 -0.165 176.285 0.165 ;
        RECT 175.96 -0.165 176.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.315 1.195 177.645 1.525 ;
        RECT 177.315 -0.165 177.645 0.165 ;
        RECT 177.32 -0.165 177.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 178.675 1.195 179.005 1.525 ;
        RECT 178.675 -0.165 179.005 0.165 ;
        RECT 178.68 -0.165 179 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.035 1.195 180.365 1.525 ;
        RECT 180.035 -0.165 180.365 0.165 ;
        RECT 180.04 -0.165 180.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 181.395 1.195 181.725 1.525 ;
        RECT 181.395 -0.165 181.725 0.165 ;
        RECT 181.4 -0.165 181.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.755 1.195 183.085 1.525 ;
        RECT 182.755 -0.165 183.085 0.165 ;
        RECT 182.76 -0.165 183.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.115 1.195 184.445 1.525 ;
        RECT 184.115 -0.165 184.445 0.165 ;
        RECT 184.12 -0.165 184.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 185.475 1.195 185.805 1.525 ;
        RECT 185.475 -0.165 185.805 0.165 ;
        RECT 185.48 -0.165 185.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.835 1.195 187.165 1.525 ;
        RECT 186.835 -0.165 187.165 0.165 ;
        RECT 186.84 -0.165 187.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.195 1.195 188.525 1.525 ;
        RECT 188.195 -0.165 188.525 0.165 ;
        RECT 188.2 -0.165 188.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.555 1.195 189.885 1.525 ;
        RECT 189.555 -0.165 189.885 0.165 ;
        RECT 189.56 -0.165 189.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.915 1.195 191.245 1.525 ;
        RECT 190.915 -0.165 191.245 0.165 ;
        RECT 190.92 -0.165 191.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.275 1.195 192.605 1.525 ;
        RECT 192.275 -0.165 192.605 0.165 ;
        RECT 192.28 -0.165 192.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 193.635 1.195 193.965 1.525 ;
        RECT 193.635 -0.165 193.965 0.165 ;
        RECT 193.64 -0.165 193.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.995 1.195 195.325 1.525 ;
        RECT 194.995 -0.165 195.325 0.165 ;
        RECT 195 -0.165 195.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 196.355 1.195 196.685 1.525 ;
        RECT 196.355 -0.165 196.685 0.165 ;
        RECT 196.36 -0.165 196.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.715 1.195 198.045 1.525 ;
        RECT 197.715 -0.165 198.045 0.165 ;
        RECT 197.72 -0.165 198.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.075 1.195 199.405 1.525 ;
        RECT 199.075 -0.165 199.405 0.165 ;
        RECT 199.08 -0.165 199.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 200.435 1.195 200.765 1.525 ;
        RECT 200.435 -0.165 200.765 0.165 ;
        RECT 200.44 -0.165 200.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.795 1.195 202.125 1.525 ;
        RECT 201.795 -0.165 202.125 0.165 ;
        RECT 201.8 -0.165 202.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.155 1.195 203.485 1.525 ;
        RECT 203.155 -0.165 203.485 0.165 ;
        RECT 203.16 -0.165 203.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 204.515 1.195 204.845 1.525 ;
        RECT 204.515 -0.165 204.845 0.165 ;
        RECT 204.52 -0.165 204.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.875 1.195 206.205 1.525 ;
        RECT 205.875 -0.165 206.205 0.165 ;
        RECT 205.88 -0.165 206.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.235 1.195 207.565 1.525 ;
        RECT 207.235 -0.165 207.565 0.165 ;
        RECT 207.24 -0.165 207.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 208.595 1.195 208.925 1.525 ;
        RECT 208.595 -0.165 208.925 0.165 ;
        RECT 208.6 -0.165 208.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.955 1.195 210.285 1.525 ;
        RECT 209.955 -0.165 210.285 0.165 ;
        RECT 209.96 -0.165 210.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 211.315 1.195 211.645 1.525 ;
        RECT 211.315 -0.165 211.645 0.165 ;
        RECT 211.32 -0.165 211.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 212.675 1.195 213.005 1.525 ;
        RECT 212.675 -0.165 213.005 0.165 ;
        RECT 212.68 -0.165 213 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.035 1.195 214.365 1.525 ;
        RECT 214.035 -0.165 214.365 0.165 ;
        RECT 214.04 -0.165 214.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 215.395 1.195 215.725 1.525 ;
        RECT 215.395 -0.165 215.725 0.165 ;
        RECT 215.4 -0.165 215.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.755 1.195 217.085 1.525 ;
        RECT 216.755 -0.165 217.085 0.165 ;
        RECT 216.76 -0.165 217.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.115 1.195 218.445 1.525 ;
        RECT 218.115 -0.165 218.445 0.165 ;
        RECT 218.12 -0.165 218.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 219.475 1.195 219.805 1.525 ;
        RECT 219.475 -0.165 219.805 0.165 ;
        RECT 219.48 -0.165 219.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.835 1.195 221.165 1.525 ;
        RECT 220.835 -0.165 221.165 0.165 ;
        RECT 220.84 -0.165 221.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.195 1.195 222.525 1.525 ;
        RECT 222.195 -0.165 222.525 0.165 ;
        RECT 222.2 -0.165 222.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 223.555 1.195 223.885 1.525 ;
        RECT 223.555 -0.165 223.885 0.165 ;
        RECT 223.56 -0.165 223.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 224.915 1.195 225.245 1.525 ;
        RECT 224.915 -0.165 225.245 0.165 ;
        RECT 224.92 -0.165 225.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.275 1.195 226.605 1.525 ;
        RECT 226.275 -0.165 226.605 0.165 ;
        RECT 226.28 -0.165 226.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 227.635 1.195 227.965 1.525 ;
        RECT 227.635 -0.165 227.965 0.165 ;
        RECT 227.64 -0.165 227.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.995 1.195 229.325 1.525 ;
        RECT 228.995 -0.165 229.325 0.165 ;
        RECT 229 -0.165 229.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 230.355 1.195 230.685 1.525 ;
        RECT 230.355 -0.165 230.685 0.165 ;
        RECT 230.36 -0.165 230.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 231.715 1.195 232.045 1.525 ;
        RECT 231.715 -0.165 232.045 0.165 ;
        RECT 231.72 -0.165 232.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.075 1.195 233.405 1.525 ;
        RECT 233.075 -0.165 233.405 0.165 ;
        RECT 233.08 -0.165 233.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 234.435 1.195 234.765 1.525 ;
        RECT 234.435 -0.165 234.765 0.165 ;
        RECT 234.44 -0.165 234.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 235.795 1.195 236.125 1.525 ;
        RECT 235.795 -0.165 236.125 0.165 ;
        RECT 235.8 -0.165 236.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 237.155 1.195 237.485 1.525 ;
        RECT 237.155 -0.165 237.485 0.165 ;
        RECT 237.16 -0.165 237.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 238.515 1.195 238.845 1.525 ;
        RECT 238.515 -0.165 238.845 0.165 ;
        RECT 238.52 -0.165 238.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.875 1.195 240.205 1.525 ;
        RECT 239.875 -0.165 240.205 0.165 ;
        RECT 239.88 -0.165 240.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 241.235 1.195 241.565 1.525 ;
        RECT 241.235 -0.165 241.565 0.165 ;
        RECT 241.24 -0.165 241.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 242.595 1.195 242.925 1.525 ;
        RECT 242.595 -0.165 242.925 0.165 ;
        RECT 242.6 -0.165 242.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 243.955 1.195 244.285 1.525 ;
        RECT 243.955 -0.165 244.285 0.165 ;
        RECT 243.96 -0.165 244.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 245.315 1.195 245.645 1.525 ;
        RECT 245.315 -0.165 245.645 0.165 ;
        RECT 245.32 -0.165 245.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 246.675 1.195 247.005 1.525 ;
        RECT 246.675 -0.165 247.005 0.165 ;
        RECT 246.68 -0.165 247 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.035 1.195 248.365 1.525 ;
        RECT 248.035 -0.165 248.365 0.165 ;
        RECT 248.04 -0.165 248.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 249.395 1.195 249.725 1.525 ;
        RECT 249.395 -0.165 249.725 0.165 ;
        RECT 249.4 -0.165 249.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.755 1.195 251.085 1.525 ;
        RECT 250.755 -0.165 251.085 0.165 ;
        RECT 250.76 -0.165 251.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.115 1.195 252.445 1.525 ;
        RECT 252.115 -0.165 252.445 0.165 ;
        RECT 252.12 -0.165 252.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 253.475 1.195 253.805 1.525 ;
        RECT 253.475 -0.165 253.805 0.165 ;
        RECT 253.48 -0.165 253.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 254.835 1.195 255.165 1.525 ;
        RECT 254.835 -0.165 255.165 0.165 ;
        RECT 254.84 -0.165 255.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 256.195 1.195 256.525 1.525 ;
        RECT 256.195 -0.165 256.525 0.165 ;
        RECT 256.2 -0.165 256.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 257.555 1.195 257.885 1.525 ;
        RECT 257.555 -0.165 257.885 0.165 ;
        RECT 257.56 -0.165 257.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.915 1.195 259.245 1.525 ;
        RECT 258.915 -0.165 259.245 0.165 ;
        RECT 258.92 -0.165 259.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.275 1.195 260.605 1.525 ;
        RECT 260.275 -0.165 260.605 0.165 ;
        RECT 260.28 -0.165 260.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 261.635 1.195 261.965 1.525 ;
        RECT 261.635 -0.165 261.965 0.165 ;
        RECT 261.64 -0.165 261.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.995 1.195 263.325 1.525 ;
        RECT 262.995 -0.165 263.325 0.165 ;
        RECT 263 -0.165 263.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 264.355 1.195 264.685 1.525 ;
        RECT 264.355 -0.165 264.685 0.165 ;
        RECT 264.36 -0.165 264.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 265.715 1.195 266.045 1.525 ;
        RECT 265.715 -0.165 266.045 0.165 ;
        RECT 265.72 -0.165 266.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 267.075 1.195 267.405 1.525 ;
        RECT 267.075 -0.165 267.405 0.165 ;
        RECT 267.08 -0.165 267.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 268.435 1.195 268.765 1.525 ;
        RECT 268.435 -0.165 268.765 0.165 ;
        RECT 268.44 -0.165 268.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.795 1.195 270.125 1.525 ;
        RECT 269.795 -0.165 270.125 0.165 ;
        RECT 269.8 -0.165 270.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.155 1.195 271.485 1.525 ;
        RECT 271.155 -0.165 271.485 0.165 ;
        RECT 271.16 -0.165 271.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 272.515 1.195 272.845 1.525 ;
        RECT 272.515 -0.165 272.845 0.165 ;
        RECT 272.52 -0.165 272.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.875 1.195 274.205 1.525 ;
        RECT 273.875 -0.165 274.205 0.165 ;
        RECT 273.88 -0.165 274.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.235 1.195 275.565 1.525 ;
        RECT 275.235 -0.165 275.565 0.165 ;
        RECT 275.24 -0.165 275.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 276.595 1.195 276.925 1.525 ;
        RECT 276.595 -0.165 276.925 0.165 ;
        RECT 276.6 -0.165 276.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 277.955 1.195 278.285 1.525 ;
        RECT 277.955 -0.165 278.285 0.165 ;
        RECT 277.96 -0.165 278.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.315 1.195 279.645 1.525 ;
        RECT 279.315 -0.165 279.645 0.165 ;
        RECT 279.32 -0.165 279.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 280.675 1.195 281.005 1.525 ;
        RECT 280.675 -0.165 281.005 0.165 ;
        RECT 280.68 -0.165 281 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.035 1.195 282.365 1.525 ;
        RECT 282.035 -0.165 282.365 0.165 ;
        RECT 282.04 -0.165 282.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 283.395 1.195 283.725 1.525 ;
        RECT 283.395 -0.165 283.725 0.165 ;
        RECT 283.4 -0.165 283.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 284.755 1.195 285.085 1.525 ;
        RECT 284.755 -0.165 285.085 0.165 ;
        RECT 284.76 -0.165 285.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.115 1.195 286.445 1.525 ;
        RECT 286.115 -0.165 286.445 0.165 ;
        RECT 286.12 -0.165 286.44 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 287.475 1.195 287.805 1.525 ;
        RECT 287.475 -0.165 287.805 0.165 ;
        RECT 287.48 -0.165 287.8 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.835 1.195 289.165 1.525 ;
        RECT 288.835 -0.165 289.165 0.165 ;
        RECT 288.84 -0.165 289.16 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.195 1.195 290.525 1.525 ;
        RECT 290.195 -0.165 290.525 0.165 ;
        RECT 290.2 -0.165 290.52 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 291.555 1.195 291.885 1.525 ;
        RECT 291.555 -0.165 291.885 0.165 ;
        RECT 291.56 -0.165 291.88 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.915 1.195 293.245 1.525 ;
        RECT 292.915 -0.165 293.245 0.165 ;
        RECT 292.92 -0.165 293.24 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.275 1.195 294.605 1.525 ;
        RECT 294.275 -0.165 294.605 0.165 ;
        RECT 294.28 -0.165 294.6 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 295.635 1.195 295.965 1.525 ;
        RECT 295.635 -0.165 295.965 0.165 ;
        RECT 295.64 -0.165 295.96 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 296.995 1.195 297.325 1.525 ;
        RECT 296.995 -0.165 297.325 0.165 ;
        RECT 297 -0.165 297.32 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 298.355 1.195 298.685 1.525 ;
        RECT 298.355 -0.165 298.685 0.165 ;
        RECT 298.36 -0.165 298.68 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 299.715 1.195 300.045 1.525 ;
        RECT 299.715 -0.165 300.045 0.165 ;
        RECT 299.72 -0.165 300.04 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.075 1.195 301.405 1.525 ;
        RECT 301.075 -0.165 301.405 0.165 ;
        RECT 301.08 -0.165 301.4 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 302.435 1.195 302.765 1.525 ;
        RECT 302.435 -0.165 302.765 0.165 ;
        RECT 302.44 -0.165 302.76 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.795 1.195 304.125 1.525 ;
        RECT 303.795 -0.165 304.125 0.165 ;
        RECT 303.8 -0.165 304.12 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.155 1.195 305.485 1.525 ;
        RECT 305.155 -0.165 305.485 0.165 ;
        RECT 305.16 -0.165 305.48 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 306.515 1.195 306.845 1.525 ;
        RECT 306.515 -0.165 306.845 0.165 ;
        RECT 306.52 -0.165 306.84 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.875 1.195 308.205 1.525 ;
        RECT 307.875 -0.165 308.205 0.165 ;
        RECT 307.88 -0.165 308.2 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.235 1.195 309.565 1.525 ;
        RECT 309.235 -0.165 309.565 0.165 ;
        RECT 309.24 -0.165 309.56 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 310.595 1.195 310.925 1.525 ;
        RECT 310.595 -0.165 310.925 0.165 ;
        RECT 310.6 -0.165 310.92 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 311.955 1.195 312.285 1.525 ;
        RECT 311.955 -0.165 312.285 0.165 ;
        RECT 311.96 -0.165 312.28 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.315 1.195 313.645 1.525 ;
        RECT 313.315 -0.165 313.645 0.165 ;
        RECT 313.32 -0.165 313.64 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 314.675 1.195 315.005 1.525 ;
        RECT 314.675 -0.165 315.005 0.165 ;
        RECT 314.68 -0.165 315 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 316.035 1.195 316.365 1.525 ;
        RECT 316.035 -0.165 316.365 0.165 ;
        RECT 316.04 -0.165 316.36 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 317.395 1.195 317.725 1.525 ;
        RECT 317.395 -0.165 317.725 0.165 ;
        RECT 317.4 -0.165 317.72 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.755 1.195 319.085 1.525 ;
        RECT 318.755 -0.165 319.085 0.165 ;
        RECT 318.76 -0.165 319.08 7.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 320.115 -0.165 320.445 0.165 ;
        RECT 320.12 -0.165 320.44 7.64 ;
        RECT 320.115 1.195 320.445 1.525 ;
    END
  END vss
  OBS
    LAYER met1 ;
      RECT 766.05 -2.4 766.37 9.32 ;
      RECT 762.03 -2.4 762.35 9.32 ;
      RECT 760.05 -2.4 760.37 9.32 ;
      RECT 756.03 -2.4 756.35 9.32 ;
      RECT 754.05 -2.4 754.37 9.32 ;
      RECT 750.03 -2.4 750.35 9.32 ;
      RECT 748.05 -2.4 748.37 9.32 ;
      RECT 744.03 -2.4 744.35 9.32 ;
      RECT 742.05 -2.4 742.37 9.32 ;
      RECT 738.03 -2.4 738.35 9.32 ;
      RECT 736.05 -2.4 736.37 9.32 ;
      RECT 732.03 -2.4 732.35 9.32 ;
      RECT 730.05 -2.4 730.37 9.32 ;
      RECT 726.03 -2.4 726.35 9.32 ;
      RECT 724.05 -2.4 724.37 9.32 ;
      RECT 720.03 -2.4 720.35 9.32 ;
      RECT 718.05 -2.4 718.37 9.32 ;
      RECT 714.03 -2.4 714.35 9.32 ;
      RECT 712.05 -2.4 712.37 9.32 ;
      RECT 708.03 -2.4 708.35 9.32 ;
      RECT 706.05 -2.4 706.37 9.32 ;
      RECT 702.03 -2.4 702.35 9.32 ;
      RECT 700.05 -2.4 700.37 9.32 ;
      RECT 696.03 -2.4 696.35 9.32 ;
      RECT 694.05 -2.4 694.37 9.32 ;
      RECT 690.03 -2.4 690.35 9.32 ;
      RECT 688.05 -2.4 688.37 9.32 ;
      RECT 684.03 -2.4 684.35 9.32 ;
      RECT 682.05 -2.4 682.37 9.32 ;
      RECT 678.03 -2.4 678.35 9.32 ;
      RECT 676.05 -2.4 676.37 9.32 ;
      RECT 672.03 -2.4 672.35 9.32 ;
      RECT 670.05 -2.4 670.37 9.32 ;
      RECT 666.03 -2.4 666.35 9.32 ;
      RECT 664.05 -2.4 664.37 9.32 ;
      RECT 660.03 -2.4 660.35 9.32 ;
      RECT 658.05 -2.4 658.37 9.32 ;
      RECT 654.03 -2.4 654.35 9.32 ;
      RECT 652.05 -2.4 652.37 9.32 ;
      RECT 648.03 -2.4 648.35 9.32 ;
      RECT 646.05 -2.4 646.37 9.32 ;
      RECT 642.03 -2.4 642.35 9.32 ;
      RECT 640.05 -2.4 640.37 9.32 ;
      RECT 636.03 -2.4 636.35 9.32 ;
      RECT 634.05 -2.4 634.37 9.32 ;
      RECT 630.03 -2.4 630.35 9.32 ;
      RECT 628.05 -2.4 628.37 9.32 ;
      RECT 624.03 -2.4 624.35 9.32 ;
      RECT 622.05 -2.4 622.37 9.32 ;
      RECT 618.03 -2.4 618.35 9.32 ;
      RECT 616.05 -2.4 616.37 9.32 ;
      RECT 612.03 -2.4 612.35 9.32 ;
      RECT 610.05 -2.4 610.37 9.32 ;
      RECT 606.03 -2.4 606.35 9.32 ;
      RECT 604.05 -2.4 604.37 9.32 ;
      RECT 600.03 -2.4 600.35 9.32 ;
      RECT 598.05 -2.4 598.37 9.32 ;
      RECT 594.03 -2.4 594.35 9.32 ;
      RECT 592.05 -2.4 592.37 9.32 ;
      RECT 588.03 -2.4 588.35 9.32 ;
      RECT 586.05 -2.4 586.37 9.32 ;
      RECT 582.03 -2.4 582.35 9.32 ;
      RECT 580.05 -2.4 580.37 9.32 ;
      RECT 576.03 -2.4 576.35 9.32 ;
      RECT 574.05 -2.4 574.37 9.32 ;
      RECT 570.03 -2.4 570.35 9.32 ;
      RECT 568.05 -2.4 568.37 9.32 ;
      RECT 564.03 -2.4 564.35 9.32 ;
      RECT 562.05 -2.4 562.37 9.32 ;
      RECT 558.03 -2.4 558.35 9.32 ;
      RECT 556.05 -2.4 556.37 9.32 ;
      RECT 552.03 -2.4 552.35 9.32 ;
      RECT 550.05 -2.4 550.37 9.32 ;
      RECT 546.03 -2.4 546.35 9.32 ;
      RECT 544.05 -2.4 544.37 9.32 ;
      RECT 540.03 -2.4 540.35 9.32 ;
      RECT 538.05 -2.4 538.37 9.32 ;
      RECT 534.03 -2.4 534.35 9.32 ;
      RECT 532.05 -2.4 532.37 9.32 ;
      RECT 528.03 -2.4 528.35 9.32 ;
      RECT 526.05 -2.4 526.37 9.32 ;
      RECT 522.03 -2.4 522.35 9.32 ;
      RECT 520.05 -2.4 520.37 9.32 ;
      RECT 516.03 -2.4 516.35 9.32 ;
      RECT 514.05 -2.4 514.37 9.32 ;
      RECT 510.03 -2.4 510.35 9.32 ;
      RECT 508.05 -2.4 508.37 9.32 ;
      RECT 504.03 -2.4 504.35 9.32 ;
      RECT 502.05 -2.4 502.37 9.32 ;
      RECT 498.03 -2.4 498.35 9.32 ;
      RECT 496.05 -2.4 496.37 9.32 ;
      RECT 492.03 -2.4 492.35 9.32 ;
      RECT 490.05 -2.4 490.37 9.32 ;
      RECT 486.03 -2.4 486.35 9.32 ;
      RECT 484.05 -2.4 484.37 9.32 ;
      RECT 480.03 -2.4 480.35 9.32 ;
      RECT 478.05 -2.4 478.37 9.32 ;
      RECT 474.03 -2.4 474.35 9.32 ;
      RECT 472.05 -2.4 472.37 9.32 ;
      RECT 468.03 -2.4 468.35 9.32 ;
      RECT 466.05 -2.4 466.37 9.32 ;
      RECT 462.03 -2.4 462.35 9.32 ;
      RECT 460.05 -2.4 460.37 9.32 ;
      RECT 456.03 -2.4 456.35 9.32 ;
      RECT 454.05 -2.4 454.37 9.32 ;
      RECT 450.03 -2.4 450.35 9.32 ;
      RECT 448.05 -2.4 448.37 9.32 ;
      RECT 444.03 -2.4 444.35 9.32 ;
      RECT 442.05 -2.4 442.37 9.32 ;
      RECT 438.03 -2.4 438.35 9.32 ;
      RECT 436.05 -2.4 436.37 9.32 ;
      RECT 432.03 -2.4 432.35 9.32 ;
      RECT 430.05 -2.4 430.37 9.32 ;
      RECT 426.03 -2.4 426.35 9.32 ;
      RECT 424.05 -2.4 424.37 9.32 ;
      RECT 420.03 -2.4 420.35 9.32 ;
      RECT 418.05 -2.4 418.37 9.32 ;
      RECT 414.03 -2.4 414.35 9.32 ;
      RECT 412.05 -2.4 412.37 9.32 ;
      RECT 408.03 -2.4 408.35 9.32 ;
      RECT 406.05 -2.4 406.37 9.32 ;
      RECT 402.03 -2.4 402.35 9.32 ;
      RECT 400.05 -2.4 400.37 9.32 ;
      RECT 396.03 -2.4 396.35 9.32 ;
      RECT 394.05 -2.4 394.37 9.32 ;
      RECT 390.03 -2.4 390.35 9.32 ;
      RECT 388.05 -2.4 388.37 9.32 ;
      RECT 384.03 -2.4 384.35 9.32 ;
      RECT 382.05 -2.4 382.37 9.32 ;
      RECT 378.03 -2.4 378.35 9.32 ;
      RECT 376.05 -2.4 376.37 9.32 ;
      RECT 372.03 -2.4 372.35 9.32 ;
      RECT 370.05 -2.4 370.37 9.32 ;
      RECT 366.03 -2.4 366.35 9.32 ;
      RECT 364.05 -2.4 364.37 9.32 ;
      RECT 360.03 -2.4 360.35 9.32 ;
      RECT 358.05 -2.4 358.37 9.32 ;
      RECT 354.03 -2.4 354.35 9.32 ;
      RECT 352.05 -2.4 352.37 9.32 ;
      RECT 348.03 -2.4 348.35 9.32 ;
      RECT 346.05 -2.4 346.37 9.32 ;
      RECT 342.03 -2.4 342.35 9.32 ;
      RECT 340.05 -2.4 340.37 9.32 ;
      RECT 336.03 -2.4 336.35 9.32 ;
      RECT 334.05 -2.4 334.37 9.32 ;
      RECT 330.03 -2.4 330.35 9.32 ;
      RECT 328.05 -2.4 328.37 9.32 ;
      RECT 324.03 -2.4 324.35 9.32 ;
      RECT 322.05 -2.4 322.37 9.32 ;
      RECT 318.03 -2.4 318.35 9.32 ;
      RECT 316.05 -2.4 316.37 9.32 ;
      RECT 312.03 -2.4 312.35 9.32 ;
      RECT 310.05 -2.4 310.37 9.32 ;
      RECT 306.03 -2.4 306.35 9.32 ;
      RECT 304.05 -2.4 304.37 9.32 ;
      RECT 300.03 -2.4 300.35 9.32 ;
      RECT 298.05 -2.4 298.37 9.32 ;
      RECT 294.03 -2.4 294.35 9.32 ;
      RECT 292.05 -2.4 292.37 9.32 ;
      RECT 288.03 -2.4 288.35 9.32 ;
      RECT 286.05 -2.4 286.37 9.32 ;
      RECT 282.03 -2.4 282.35 9.32 ;
      RECT 280.05 -2.4 280.37 9.32 ;
      RECT 276.03 -2.4 276.35 9.32 ;
      RECT 274.05 -2.4 274.37 9.32 ;
      RECT 270.03 -2.4 270.35 9.32 ;
      RECT 268.05 -2.4 268.37 9.32 ;
      RECT 264.03 -2.4 264.35 9.32 ;
      RECT 262.05 -2.4 262.37 9.32 ;
      RECT 258.03 -2.4 258.35 9.32 ;
      RECT 256.05 -2.4 256.37 9.32 ;
      RECT 252.03 -2.4 252.35 9.32 ;
      RECT 250.05 -2.4 250.37 9.32 ;
      RECT 246.03 -2.4 246.35 9.32 ;
      RECT 244.05 -2.4 244.37 9.32 ;
      RECT 240.03 -2.4 240.35 9.32 ;
      RECT 238.05 -2.4 238.37 9.32 ;
      RECT 234.03 -2.4 234.35 9.32 ;
      RECT 232.05 -2.4 232.37 9.32 ;
      RECT 228.03 -2.4 228.35 9.32 ;
      RECT 226.05 -2.4 226.37 9.32 ;
      RECT 222.03 -2.4 222.35 9.32 ;
      RECT 220.05 -2.4 220.37 9.32 ;
      RECT 216.03 -2.4 216.35 9.32 ;
      RECT 214.05 -2.4 214.37 9.32 ;
      RECT 210.03 -2.4 210.35 9.32 ;
      RECT 208.05 -2.4 208.37 9.32 ;
      RECT 204.03 -2.4 204.35 9.32 ;
      RECT 202.05 -2.4 202.37 9.32 ;
      RECT 198.03 -2.4 198.35 9.32 ;
      RECT 196.05 -2.4 196.37 9.32 ;
      RECT 192.03 -2.4 192.35 9.32 ;
      RECT 190.05 -2.4 190.37 9.32 ;
      RECT 186.03 -2.4 186.35 9.32 ;
      RECT 184.05 -2.4 184.37 9.32 ;
      RECT 180.03 -2.4 180.35 9.32 ;
      RECT 178.05 -2.4 178.37 9.32 ;
      RECT 174.03 -2.4 174.35 9.32 ;
      RECT 172.05 -2.4 172.37 9.32 ;
      RECT 168.03 -2.4 168.35 9.32 ;
      RECT 166.05 -2.4 166.37 9.32 ;
      RECT 162.03 -2.4 162.35 9.32 ;
      RECT 160.05 -2.4 160.37 9.32 ;
      RECT 156.03 -2.4 156.35 9.32 ;
      RECT 154.05 -2.4 154.37 9.32 ;
      RECT 150.03 -2.4 150.35 9.32 ;
      RECT 148.05 -2.4 148.37 9.32 ;
      RECT 144.03 -2.4 144.35 9.32 ;
      RECT 142.05 -2.4 142.37 9.32 ;
      RECT 138.03 -2.4 138.35 9.32 ;
      RECT 136.05 -2.4 136.37 9.32 ;
      RECT 132.03 -2.4 132.35 9.32 ;
      RECT 130.05 -2.4 130.37 9.32 ;
      RECT 126.03 -2.4 126.35 9.32 ;
      RECT 124.05 -2.4 124.37 9.32 ;
      RECT 120.03 -2.4 120.35 9.32 ;
      RECT 118.05 -2.4 118.37 9.32 ;
      RECT 114.03 -2.4 114.35 9.32 ;
      RECT 112.05 -2.4 112.37 9.32 ;
      RECT 108.03 -2.4 108.35 9.32 ;
      RECT 106.05 -2.4 106.37 9.32 ;
      RECT 102.03 -2.4 102.35 9.32 ;
      RECT 100.05 -2.4 100.37 9.32 ;
      RECT 96.03 -2.4 96.35 9.32 ;
      RECT 94.05 -2.4 94.37 9.32 ;
      RECT 90.03 -2.4 90.35 9.32 ;
      RECT 88.05 -2.4 88.37 9.32 ;
      RECT 84.03 -2.4 84.35 9.32 ;
      RECT 82.05 -2.4 82.37 9.32 ;
      RECT 78.03 -2.4 78.35 9.32 ;
      RECT 76.05 -2.4 76.37 9.32 ;
      RECT 72.03 -2.4 72.35 9.32 ;
      RECT 70.05 -2.4 70.37 9.32 ;
      RECT 66.03 -2.4 66.35 9.32 ;
      RECT 64.05 -2.4 64.37 9.32 ;
      RECT 60.03 -2.4 60.35 9.32 ;
      RECT 58.05 -2.4 58.37 9.32 ;
      RECT 54.03 -2.4 54.35 9.32 ;
      RECT 52.05 -2.4 52.37 9.32 ;
      RECT 48.03 -2.4 48.35 9.32 ;
      RECT 46.05 -2.4 46.37 9.32 ;
      RECT 42.03 -2.4 42.35 9.32 ;
      RECT 40.05 -2.4 40.37 9.32 ;
      RECT 36.03 -2.4 36.35 9.32 ;
      RECT 34.05 -2.4 34.37 9.32 ;
      RECT 30.03 -2.4 30.35 9.32 ;
      RECT 28.05 -2.4 28.37 9.32 ;
      RECT 24.03 -2.4 24.35 9.32 ;
      RECT 22.05 -2.4 22.37 9.32 ;
      RECT 18.03 -2.4 18.35 9.32 ;
      RECT 16.05 -2.4 16.37 9.32 ;
      RECT 12.03 -2.4 12.35 9.32 ;
      RECT 10.05 -2.4 10.37 9.32 ;
      RECT 6.03 -2.4 6.35 9.32 ;
      RECT 4.05 -2.4 4.37 9.32 ;
      RECT 1.52 -2.4 1.84 9.32 ;
      RECT 0.03 -2.4 0.35 9.32 ;
      RECT -1.47 -2.4 -1.15 9.32 ;
    LAYER met1 SPACING 0.14 ;
      RECT 766.67 -3 769.945 9.92 ;
      RECT 762.65 -3 765.75 9.92 ;
      RECT 760.67 -3 761.73 9.92 ;
      RECT 756.65 -3 759.75 9.92 ;
      RECT 754.67 -3 755.73 9.92 ;
      RECT 750.65 -3 753.75 9.92 ;
      RECT 748.67 -3 749.73 9.92 ;
      RECT 744.65 -3 747.75 9.92 ;
      RECT 742.67 -3 743.73 9.92 ;
      RECT 738.65 -3 741.75 9.92 ;
      RECT 736.67 -3 737.73 9.92 ;
      RECT 732.65 -3 735.75 9.92 ;
      RECT 730.67 -3 731.73 9.92 ;
      RECT 726.65 -3 729.75 9.92 ;
      RECT 724.67 -3 725.73 9.92 ;
      RECT 720.65 -3 723.75 9.92 ;
      RECT 718.67 -3 719.73 9.92 ;
      RECT 714.65 -3 717.75 9.92 ;
      RECT 712.67 -3 713.73 9.92 ;
      RECT 708.65 -3 711.75 9.92 ;
      RECT 706.67 -3 707.73 9.92 ;
      RECT 702.65 -3 705.75 9.92 ;
      RECT 700.67 -3 701.73 9.92 ;
      RECT 696.65 -3 699.75 9.92 ;
      RECT 694.67 -3 695.73 9.92 ;
      RECT 690.65 -3 693.75 9.92 ;
      RECT 688.67 -3 689.73 9.92 ;
      RECT 684.65 -3 687.75 9.92 ;
      RECT 682.67 -3 683.73 9.92 ;
      RECT 678.65 -3 681.75 9.92 ;
      RECT 676.67 -3 677.73 9.92 ;
      RECT 672.65 -3 675.75 9.92 ;
      RECT 670.67 -3 671.73 9.92 ;
      RECT 666.65 -3 669.75 9.92 ;
      RECT 664.67 -3 665.73 9.92 ;
      RECT 660.65 -3 663.75 9.92 ;
      RECT 658.67 -3 659.73 9.92 ;
      RECT 654.65 -3 657.75 9.92 ;
      RECT 652.67 -3 653.73 9.92 ;
      RECT 648.65 -3 651.75 9.92 ;
      RECT 646.67 -3 647.73 9.92 ;
      RECT 642.65 -3 645.75 9.92 ;
      RECT 640.67 -3 641.73 9.92 ;
      RECT 636.65 -3 639.75 9.92 ;
      RECT 634.67 -3 635.73 9.92 ;
      RECT 630.65 -3 633.75 9.92 ;
      RECT 628.67 -3 629.73 9.92 ;
      RECT 624.65 -3 627.75 9.92 ;
      RECT 622.67 -3 623.73 9.92 ;
      RECT 618.65 -3 621.75 9.92 ;
      RECT 616.67 -3 617.73 9.92 ;
      RECT 612.65 -3 615.75 9.92 ;
      RECT 610.67 -3 611.73 9.92 ;
      RECT 606.65 -3 609.75 9.92 ;
      RECT 604.67 -3 605.73 9.92 ;
      RECT 600.65 -3 603.75 9.92 ;
      RECT 598.67 -3 599.73 9.92 ;
      RECT 594.65 -3 597.75 9.92 ;
      RECT 592.67 -3 593.73 9.92 ;
      RECT 588.65 -3 591.75 9.92 ;
      RECT 586.67 -3 587.73 9.92 ;
      RECT 582.65 -3 585.75 9.92 ;
      RECT 580.67 -3 581.73 9.92 ;
      RECT 576.65 -3 579.75 9.92 ;
      RECT 574.67 -3 575.73 9.92 ;
      RECT 570.65 -3 573.75 9.92 ;
      RECT 568.67 -3 569.73 9.92 ;
      RECT 564.65 -3 567.75 9.92 ;
      RECT 562.67 -3 563.73 9.92 ;
      RECT 558.65 -3 561.75 9.92 ;
      RECT 556.67 -3 557.73 9.92 ;
      RECT 552.65 -3 555.75 9.92 ;
      RECT 550.67 -3 551.73 9.92 ;
      RECT 546.65 -3 549.75 9.92 ;
      RECT 544.67 -3 545.73 9.92 ;
      RECT 540.65 -3 543.75 9.92 ;
      RECT 538.67 -3 539.73 9.92 ;
      RECT 534.65 -3 537.75 9.92 ;
      RECT 532.67 -3 533.73 9.92 ;
      RECT 528.65 -3 531.75 9.92 ;
      RECT 526.67 -3 527.73 9.92 ;
      RECT 522.65 -3 525.75 9.92 ;
      RECT 520.67 -3 521.73 9.92 ;
      RECT 516.65 -3 519.75 9.92 ;
      RECT 514.67 -3 515.73 9.92 ;
      RECT 510.65 -3 513.75 9.92 ;
      RECT 508.67 -3 509.73 9.92 ;
      RECT 504.65 -3 507.75 9.92 ;
      RECT 502.67 -3 503.73 9.92 ;
      RECT 498.65 -3 501.75 9.92 ;
      RECT 496.67 -3 497.73 9.92 ;
      RECT 492.65 -3 495.75 9.92 ;
      RECT 490.67 -3 491.73 9.92 ;
      RECT 486.65 -3 489.75 9.92 ;
      RECT 484.67 -3 485.73 9.92 ;
      RECT 480.65 -3 483.75 9.92 ;
      RECT 478.67 -3 479.73 9.92 ;
      RECT 474.65 -3 477.75 9.92 ;
      RECT 472.67 -3 473.73 9.92 ;
      RECT 468.65 -3 471.75 9.92 ;
      RECT 466.67 -3 467.73 9.92 ;
      RECT 462.65 -3 465.75 9.92 ;
      RECT 460.67 -3 461.73 9.92 ;
      RECT 456.65 -3 459.75 9.92 ;
      RECT 454.67 -3 455.73 9.92 ;
      RECT 450.65 -3 453.75 9.92 ;
      RECT 448.67 -3 449.73 9.92 ;
      RECT 444.65 -3 447.75 9.92 ;
      RECT 442.67 -3 443.73 9.92 ;
      RECT 438.65 -3 441.75 9.92 ;
      RECT 436.67 -3 437.73 9.92 ;
      RECT 432.65 -3 435.75 9.92 ;
      RECT 430.67 -3 431.73 9.92 ;
      RECT 426.65 -3 429.75 9.92 ;
      RECT 424.67 -3 425.73 9.92 ;
      RECT 420.65 -3 423.75 9.92 ;
      RECT 418.67 -3 419.73 9.92 ;
      RECT 414.65 -3 417.75 9.92 ;
      RECT 412.67 -3 413.73 9.92 ;
      RECT 408.65 -3 411.75 9.92 ;
      RECT 406.67 -3 407.73 9.92 ;
      RECT 402.65 -3 405.75 9.92 ;
      RECT 400.67 -3 401.73 9.92 ;
      RECT 396.65 -3 399.75 9.92 ;
      RECT 394.67 -3 395.73 9.92 ;
      RECT 390.65 -3 393.75 9.92 ;
      RECT 388.67 -3 389.73 9.92 ;
      RECT 384.65 -3 387.75 9.92 ;
      RECT 382.67 -3 383.73 9.92 ;
      RECT 378.65 -3 381.75 9.92 ;
      RECT 376.67 -3 377.73 9.92 ;
      RECT 372.65 -3 375.75 9.92 ;
      RECT 370.67 -3 371.73 9.92 ;
      RECT 366.65 -3 369.75 9.92 ;
      RECT 364.67 -3 365.73 9.92 ;
      RECT 360.65 -3 363.75 9.92 ;
      RECT 358.67 -3 359.73 9.92 ;
      RECT 354.65 -3 357.75 9.92 ;
      RECT 352.67 -3 353.73 9.92 ;
      RECT 348.65 -3 351.75 9.92 ;
      RECT 346.67 -3 347.73 9.92 ;
      RECT 342.65 -3 345.75 9.92 ;
      RECT 340.67 -3 341.73 9.92 ;
      RECT 336.65 -3 339.75 9.92 ;
      RECT 334.67 -3 335.73 9.92 ;
      RECT 330.65 -3 333.75 9.92 ;
      RECT 328.67 -3 329.73 9.92 ;
      RECT 324.65 -3 327.75 9.92 ;
      RECT 322.67 -3 323.73 9.92 ;
      RECT 318.65 -3 321.75 9.92 ;
      RECT 316.67 -3 317.73 9.92 ;
      RECT 312.65 -3 315.75 9.92 ;
      RECT 310.67 -3 311.73 9.92 ;
      RECT 306.65 -3 309.75 9.92 ;
      RECT 304.67 -3 305.73 9.92 ;
      RECT 300.65 -3 303.75 9.92 ;
      RECT 298.67 -3 299.73 9.92 ;
      RECT 294.65 -3 297.75 9.92 ;
      RECT 292.67 -3 293.73 9.92 ;
      RECT 288.65 -3 291.75 9.92 ;
      RECT 286.67 -3 287.73 9.92 ;
      RECT 282.65 -3 285.75 9.92 ;
      RECT 280.67 -3 281.73 9.92 ;
      RECT 276.65 -3 279.75 9.92 ;
      RECT 274.67 -3 275.73 9.92 ;
      RECT 270.65 -3 273.75 9.92 ;
      RECT 268.67 -3 269.73 9.92 ;
      RECT 264.65 -3 267.75 9.92 ;
      RECT 262.67 -3 263.73 9.92 ;
      RECT 258.65 -3 261.75 9.92 ;
      RECT 256.67 -3 257.73 9.92 ;
      RECT 252.65 -3 255.75 9.92 ;
      RECT 250.67 -3 251.73 9.92 ;
      RECT 246.65 -3 249.75 9.92 ;
      RECT 244.67 -3 245.73 9.92 ;
      RECT 240.65 -3 243.75 9.92 ;
      RECT 238.67 -3 239.73 9.92 ;
      RECT 234.65 -3 237.75 9.92 ;
      RECT 232.67 -3 233.73 9.92 ;
      RECT 228.65 -3 231.75 9.92 ;
      RECT 226.67 -3 227.73 9.92 ;
      RECT 222.65 -3 225.75 9.92 ;
      RECT 220.67 -3 221.73 9.92 ;
      RECT 216.65 -3 219.75 9.92 ;
      RECT 214.67 -3 215.73 9.92 ;
      RECT 210.65 -3 213.75 9.92 ;
      RECT 208.67 -3 209.73 9.92 ;
      RECT 204.65 -3 207.75 9.92 ;
      RECT 202.67 -3 203.73 9.92 ;
      RECT 198.65 -3 201.75 9.92 ;
      RECT 196.67 -3 197.73 9.92 ;
      RECT 192.65 -3 195.75 9.92 ;
      RECT 190.67 -3 191.73 9.92 ;
      RECT 186.65 -3 189.75 9.92 ;
      RECT 184.67 -3 185.73 9.92 ;
      RECT 180.65 -3 183.75 9.92 ;
      RECT 178.67 -3 179.73 9.92 ;
      RECT 174.65 -3 177.75 9.92 ;
      RECT 172.67 -3 173.73 9.92 ;
      RECT 168.65 -3 171.75 9.92 ;
      RECT 166.67 -3 167.73 9.92 ;
      RECT 162.65 -3 165.75 9.92 ;
      RECT 160.67 -3 161.73 9.92 ;
      RECT 156.65 -3 159.75 9.92 ;
      RECT 154.67 -3 155.73 9.92 ;
      RECT 150.65 -3 153.75 9.92 ;
      RECT 148.67 -3 149.73 9.92 ;
      RECT 144.65 -3 147.75 9.92 ;
      RECT 142.67 -3 143.73 9.92 ;
      RECT 138.65 -3 141.75 9.92 ;
      RECT 136.67 -3 137.73 9.92 ;
      RECT 132.65 -3 135.75 9.92 ;
      RECT 130.67 -3 131.73 9.92 ;
      RECT 126.65 -3 129.75 9.92 ;
      RECT 124.67 -3 125.73 9.92 ;
      RECT 120.65 -3 123.75 9.92 ;
      RECT 118.67 -3 119.73 9.92 ;
      RECT 114.65 -3 117.75 9.92 ;
      RECT 112.67 -3 113.73 9.92 ;
      RECT 108.65 -3 111.75 9.92 ;
      RECT 106.67 -3 107.73 9.92 ;
      RECT 102.65 -3 105.75 9.92 ;
      RECT 100.67 -3 101.73 9.92 ;
      RECT 96.65 -3 99.75 9.92 ;
      RECT 94.67 -3 95.73 9.92 ;
      RECT 90.65 -3 93.75 9.92 ;
      RECT 88.67 -3 89.73 9.92 ;
      RECT 84.65 -3 87.75 9.92 ;
      RECT 82.67 -3 83.73 9.92 ;
      RECT 78.65 -3 81.75 9.92 ;
      RECT 76.67 -3 77.73 9.92 ;
      RECT 72.65 -3 75.75 9.92 ;
      RECT 70.67 -3 71.73 9.92 ;
      RECT 66.65 -3 69.75 9.92 ;
      RECT 64.67 -3 65.73 9.92 ;
      RECT 60.65 -3 63.75 9.92 ;
      RECT 58.67 -3 59.73 9.92 ;
      RECT 54.65 -3 57.75 9.92 ;
      RECT 52.67 -3 53.73 9.92 ;
      RECT 48.65 -3 51.75 9.92 ;
      RECT 46.67 -3 47.73 9.92 ;
      RECT 42.65 -3 45.75 9.92 ;
      RECT 40.67 -3 41.73 9.92 ;
      RECT 36.65 -3 39.75 9.92 ;
      RECT 34.67 -3 35.73 9.92 ;
      RECT 30.65 -3 33.75 9.92 ;
      RECT 28.67 -3 29.73 9.92 ;
      RECT 24.65 -3 27.75 9.92 ;
      RECT 22.67 -3 23.73 9.92 ;
      RECT 18.65 -3 21.75 9.92 ;
      RECT 16.67 -3 17.73 9.92 ;
      RECT 12.65 -3 15.75 9.92 ;
      RECT 10.67 -3 11.73 9.92 ;
      RECT 6.65 -3 9.75 9.92 ;
      RECT 4.67 -3 5.73 9.92 ;
      RECT 2.14 -3 3.75 9.92 ;
      RECT 0.65 -3 1.22 9.92 ;
      RECT -0.85 -3 -0.27 9.92 ;
      RECT -2.88 -3 -1.77 9.92 ;
      RECT -2.88 -2.38 769.945 9.3 ;
    LAYER met2 ;
      RECT 769.575 -0.82 769.945 -0.54 ;
      RECT 769.575 0.54 769.945 0.82 ;
      RECT 769.575 1.9 769.945 2.18 ;
      RECT 769.575 3.26 769.945 3.54 ;
      RECT 769.575 4.62 769.945 4.9 ;
      RECT 769.575 5.98 769.945 6.26 ;
      RECT -2.88 -0.16 769.24 0.16 ;
      RECT -2.88 0.52 769.24 0.84 ;
      RECT -2.88 1.2 769.24 1.52 ;
      RECT -2.88 1.88 769.24 2.2 ;
      RECT -2.88 2.56 769.24 2.88 ;
      RECT -2.88 7.32 769.24 7.64 ;
      RECT -2.88 3.24 6.96 3.56 ;
      RECT -2.88 5.28 3.56 5.6 ;
      RECT -2.88 3.92 0.84 4.24 ;
      RECT -2.88 4.6 0.84 4.92 ;
      RECT -2.88 5.96 -0.52 6.28 ;
      RECT -2.88 6.64 -0.52 6.96 ;
    LAYER met2 SPACING 0.14 ;
      RECT 766.67 -3 769.945 9.92 ;
      RECT 762.65 -3 765.75 9.92 ;
      RECT 760.67 -3 761.73 9.92 ;
      RECT 756.65 -3 759.75 9.92 ;
      RECT 754.67 -3 755.73 9.92 ;
      RECT 750.65 -3 753.75 9.92 ;
      RECT 748.67 -3 749.73 9.92 ;
      RECT 744.65 -3 747.75 9.92 ;
      RECT 742.67 -3 743.73 9.92 ;
      RECT 738.65 -3 741.75 9.92 ;
      RECT 736.67 -3 737.73 9.92 ;
      RECT 732.65 -3 735.75 9.92 ;
      RECT 730.67 -3 731.73 9.92 ;
      RECT 726.65 -3 729.75 9.92 ;
      RECT 724.67 -3 725.73 9.92 ;
      RECT 720.65 -3 723.75 9.92 ;
      RECT 718.67 -3 719.73 9.92 ;
      RECT 714.65 -3 717.75 9.92 ;
      RECT 712.67 -3 713.73 9.92 ;
      RECT 708.65 -3 711.75 9.92 ;
      RECT 706.67 -3 707.73 9.92 ;
      RECT 702.65 -3 705.75 9.92 ;
      RECT 700.67 -3 701.73 9.92 ;
      RECT 696.65 -3 699.75 9.92 ;
      RECT 694.67 -3 695.73 9.92 ;
      RECT 690.65 -3 693.75 9.92 ;
      RECT 688.67 -3 689.73 9.92 ;
      RECT 684.65 -3 687.75 9.92 ;
      RECT 682.67 -3 683.73 9.92 ;
      RECT 678.65 -3 681.75 9.92 ;
      RECT 676.67 -3 677.73 9.92 ;
      RECT 672.65 -3 675.75 9.92 ;
      RECT 670.67 -3 671.73 9.92 ;
      RECT 666.65 -3 669.75 9.92 ;
      RECT 664.67 -3 665.73 9.92 ;
      RECT 660.65 -3 663.75 9.92 ;
      RECT 658.67 -3 659.73 9.92 ;
      RECT 654.65 -3 657.75 9.92 ;
      RECT 652.67 -3 653.73 9.92 ;
      RECT 648.65 -3 651.75 9.92 ;
      RECT 646.67 -3 647.73 9.92 ;
      RECT 642.65 -3 645.75 9.92 ;
      RECT 640.67 -3 641.73 9.92 ;
      RECT 636.65 -3 639.75 9.92 ;
      RECT 634.67 -3 635.73 9.92 ;
      RECT 630.65 -3 633.75 9.92 ;
      RECT 628.67 -3 629.73 9.92 ;
      RECT 624.65 -3 627.75 9.92 ;
      RECT 622.67 -3 623.73 9.92 ;
      RECT 618.65 -3 621.75 9.92 ;
      RECT 616.67 -3 617.73 9.92 ;
      RECT 612.65 -3 615.75 9.92 ;
      RECT 610.67 -3 611.73 9.92 ;
      RECT 606.65 -3 609.75 9.92 ;
      RECT 604.67 -3 605.73 9.92 ;
      RECT 600.65 -3 603.75 9.92 ;
      RECT 598.67 -3 599.73 9.92 ;
      RECT 594.65 -3 597.75 9.92 ;
      RECT 592.67 -3 593.73 9.92 ;
      RECT 588.65 -3 591.75 9.92 ;
      RECT 586.67 -3 587.73 9.92 ;
      RECT 582.65 -3 585.75 9.92 ;
      RECT 580.67 -3 581.73 9.92 ;
      RECT 576.65 -3 579.75 9.92 ;
      RECT 574.67 -3 575.73 9.92 ;
      RECT 570.65 -3 573.75 9.92 ;
      RECT 568.67 -3 569.73 9.92 ;
      RECT 564.65 -3 567.75 9.92 ;
      RECT 562.67 -3 563.73 9.92 ;
      RECT 558.65 -3 561.75 9.92 ;
      RECT 556.67 -3 557.73 9.92 ;
      RECT 552.65 -3 555.75 9.92 ;
      RECT 550.67 -3 551.73 9.92 ;
      RECT 546.65 -3 549.75 9.92 ;
      RECT 544.67 -3 545.73 9.92 ;
      RECT 540.65 -3 543.75 9.92 ;
      RECT 538.67 -3 539.73 9.92 ;
      RECT 534.65 -3 537.75 9.92 ;
      RECT 532.67 -3 533.73 9.92 ;
      RECT 528.65 -3 531.75 9.92 ;
      RECT 526.67 -3 527.73 9.92 ;
      RECT 522.65 -3 525.75 9.92 ;
      RECT 520.67 -3 521.73 9.92 ;
      RECT 516.65 -3 519.75 9.92 ;
      RECT 514.67 -3 515.73 9.92 ;
      RECT 510.65 -3 513.75 9.92 ;
      RECT 508.67 -3 509.73 9.92 ;
      RECT 504.65 -3 507.75 9.92 ;
      RECT 502.67 -3 503.73 9.92 ;
      RECT 498.65 -3 501.75 9.92 ;
      RECT 496.67 -3 497.73 9.92 ;
      RECT 492.65 -3 495.75 9.92 ;
      RECT 490.67 -3 491.73 9.92 ;
      RECT 486.65 -3 489.75 9.92 ;
      RECT 484.67 -3 485.73 9.92 ;
      RECT 480.65 -3 483.75 9.92 ;
      RECT 478.67 -3 479.73 9.92 ;
      RECT 474.65 -3 477.75 9.92 ;
      RECT 472.67 -3 473.73 9.92 ;
      RECT 468.65 -3 471.75 9.92 ;
      RECT 466.67 -3 467.73 9.92 ;
      RECT 462.65 -3 465.75 9.92 ;
      RECT 460.67 -3 461.73 9.92 ;
      RECT 456.65 -3 459.75 9.92 ;
      RECT 454.67 -3 455.73 9.92 ;
      RECT 450.65 -3 453.75 9.92 ;
      RECT 448.67 -3 449.73 9.92 ;
      RECT 444.65 -3 447.75 9.92 ;
      RECT 442.67 -3 443.73 9.92 ;
      RECT 438.65 -3 441.75 9.92 ;
      RECT 436.67 -3 437.73 9.92 ;
      RECT 432.65 -3 435.75 9.92 ;
      RECT 430.67 -3 431.73 9.92 ;
      RECT 426.65 -3 429.75 9.92 ;
      RECT 424.67 -3 425.73 9.92 ;
      RECT 420.65 -3 423.75 9.92 ;
      RECT 418.67 -3 419.73 9.92 ;
      RECT 414.65 -3 417.75 9.92 ;
      RECT 412.67 -3 413.73 9.92 ;
      RECT 408.65 -3 411.75 9.92 ;
      RECT 406.67 -3 407.73 9.92 ;
      RECT 402.65 -3 405.75 9.92 ;
      RECT 400.67 -3 401.73 9.92 ;
      RECT 396.65 -3 399.75 9.92 ;
      RECT 394.67 -3 395.73 9.92 ;
      RECT 390.65 -3 393.75 9.92 ;
      RECT 388.67 -3 389.73 9.92 ;
      RECT 384.65 -3 387.75 9.92 ;
      RECT 382.67 -3 383.73 9.92 ;
      RECT 378.65 -3 381.75 9.92 ;
      RECT 376.67 -3 377.73 9.92 ;
      RECT 372.65 -3 375.75 9.92 ;
      RECT 370.67 -3 371.73 9.92 ;
      RECT 366.65 -3 369.75 9.92 ;
      RECT 364.67 -3 365.73 9.92 ;
      RECT 360.65 -3 363.75 9.92 ;
      RECT 358.67 -3 359.73 9.92 ;
      RECT 354.65 -3 357.75 9.92 ;
      RECT 352.67 -3 353.73 9.92 ;
      RECT 348.65 -3 351.75 9.92 ;
      RECT 346.67 -3 347.73 9.92 ;
      RECT 342.65 -3 345.75 9.92 ;
      RECT 340.67 -3 341.73 9.92 ;
      RECT 336.65 -3 339.75 9.92 ;
      RECT 334.67 -3 335.73 9.92 ;
      RECT 330.65 -3 333.75 9.92 ;
      RECT 328.67 -3 329.73 9.92 ;
      RECT 324.65 -3 327.75 9.92 ;
      RECT 322.67 -3 323.73 9.92 ;
      RECT 318.65 -3 321.75 9.92 ;
      RECT 316.67 -3 317.73 9.92 ;
      RECT 312.65 -3 315.75 9.92 ;
      RECT 310.67 -3 311.73 9.92 ;
      RECT 306.65 -3 309.75 9.92 ;
      RECT 304.67 -3 305.73 9.92 ;
      RECT 300.65 -3 303.75 9.92 ;
      RECT 298.67 -3 299.73 9.92 ;
      RECT 294.65 -3 297.75 9.92 ;
      RECT 292.67 -3 293.73 9.92 ;
      RECT 288.65 -3 291.75 9.92 ;
      RECT 286.67 -3 287.73 9.92 ;
      RECT 282.65 -3 285.75 9.92 ;
      RECT 280.67 -3 281.73 9.92 ;
      RECT 276.65 -3 279.75 9.92 ;
      RECT 274.67 -3 275.73 9.92 ;
      RECT 270.65 -3 273.75 9.92 ;
      RECT 268.67 -3 269.73 9.92 ;
      RECT 264.65 -3 267.75 9.92 ;
      RECT 262.67 -3 263.73 9.92 ;
      RECT 258.65 -3 261.75 9.92 ;
      RECT 256.67 -3 257.73 9.92 ;
      RECT 252.65 -3 255.75 9.92 ;
      RECT 250.67 -3 251.73 9.92 ;
      RECT 246.65 -3 249.75 9.92 ;
      RECT 244.67 -3 245.73 9.92 ;
      RECT 240.65 -3 243.75 9.92 ;
      RECT 238.67 -3 239.73 9.92 ;
      RECT 234.65 -3 237.75 9.92 ;
      RECT 232.67 -3 233.73 9.92 ;
      RECT 228.65 -3 231.75 9.92 ;
      RECT 226.67 -3 227.73 9.92 ;
      RECT 222.65 -3 225.75 9.92 ;
      RECT 220.67 -3 221.73 9.92 ;
      RECT 216.65 -3 219.75 9.92 ;
      RECT 214.67 -3 215.73 9.92 ;
      RECT 210.65 -3 213.75 9.92 ;
      RECT 208.67 -3 209.73 9.92 ;
      RECT 204.65 -3 207.75 9.92 ;
      RECT 202.67 -3 203.73 9.92 ;
      RECT 198.65 -3 201.75 9.92 ;
      RECT 196.67 -3 197.73 9.92 ;
      RECT 192.65 -3 195.75 9.92 ;
      RECT 190.67 -3 191.73 9.92 ;
      RECT 186.65 -3 189.75 9.92 ;
      RECT 184.67 -3 185.73 9.92 ;
      RECT 180.65 -3 183.75 9.92 ;
      RECT 178.67 -3 179.73 9.92 ;
      RECT 174.65 -3 177.75 9.92 ;
      RECT 172.67 -3 173.73 9.92 ;
      RECT 168.65 -3 171.75 9.92 ;
      RECT 166.67 -3 167.73 9.92 ;
      RECT 162.65 -3 165.75 9.92 ;
      RECT 160.67 -3 161.73 9.92 ;
      RECT 156.65 -3 159.75 9.92 ;
      RECT 154.67 -3 155.73 9.92 ;
      RECT 150.65 -3 153.75 9.92 ;
      RECT 148.67 -3 149.73 9.92 ;
      RECT 144.65 -3 147.75 9.92 ;
      RECT 142.67 -3 143.73 9.92 ;
      RECT 138.65 -3 141.75 9.92 ;
      RECT 136.67 -3 137.73 9.92 ;
      RECT 132.65 -3 135.75 9.92 ;
      RECT 130.67 -3 131.73 9.92 ;
      RECT 126.65 -3 129.75 9.92 ;
      RECT 124.67 -3 125.73 9.92 ;
      RECT 120.65 -3 123.75 9.92 ;
      RECT 118.67 -3 119.73 9.92 ;
      RECT 114.65 -3 117.75 9.92 ;
      RECT 112.67 -3 113.73 9.92 ;
      RECT 108.65 -3 111.75 9.92 ;
      RECT 106.67 -3 107.73 9.92 ;
      RECT 102.65 -3 105.75 9.92 ;
      RECT 100.67 -3 101.73 9.92 ;
      RECT 96.65 -3 99.75 9.92 ;
      RECT 94.67 -3 95.73 9.92 ;
      RECT 90.65 -3 93.75 9.92 ;
      RECT 88.67 -3 89.73 9.92 ;
      RECT 84.65 -3 87.75 9.92 ;
      RECT 82.67 -3 83.73 9.92 ;
      RECT 78.65 -3 81.75 9.92 ;
      RECT 76.67 -3 77.73 9.92 ;
      RECT 72.65 -3 75.75 9.92 ;
      RECT 70.67 -3 71.73 9.92 ;
      RECT 66.65 -3 69.75 9.92 ;
      RECT 64.67 -3 65.73 9.92 ;
      RECT 60.65 -3 63.75 9.92 ;
      RECT 58.67 -3 59.73 9.92 ;
      RECT 54.65 -3 57.75 9.92 ;
      RECT 52.67 -3 53.73 9.92 ;
      RECT 48.65 -3 51.75 9.92 ;
      RECT 46.67 -3 47.73 9.92 ;
      RECT 42.65 -3 45.75 9.92 ;
      RECT 40.67 -3 41.73 9.92 ;
      RECT 36.65 -3 39.75 9.92 ;
      RECT 34.67 -3 35.73 9.92 ;
      RECT 30.65 -3 33.75 9.92 ;
      RECT 28.67 -3 29.73 9.92 ;
      RECT 24.65 -3 27.75 9.92 ;
      RECT 22.67 -3 23.73 9.92 ;
      RECT 18.65 -3 21.75 9.92 ;
      RECT 16.67 -3 17.73 9.92 ;
      RECT 12.65 -3 15.75 9.92 ;
      RECT 10.67 -3 11.73 9.92 ;
      RECT 6.65 -3 9.75 9.92 ;
      RECT 4.67 -3 5.73 9.92 ;
      RECT 2.14 -3 3.75 9.92 ;
      RECT 0.65 -3 1.22 9.92 ;
      RECT -0.85 -3 -0.27 9.92 ;
      RECT -2.88 -3 -1.77 9.92 ;
      RECT -2.88 -2.38 769.945 9.3 ;
    LAYER met3 SPACING 0.3 ;
      RECT 769.595 -0.845 769.925 -0.515 ;
      RECT 769.595 0.515 769.925 0.845 ;
      RECT 769.595 1.875 769.925 2.205 ;
      RECT 769.595 3.235 769.925 3.565 ;
      RECT 769.595 4.595 769.925 4.925 ;
      RECT 769.595 5.955 769.925 6.285 ;
      RECT 768.915 -1.525 769.245 -1.195 ;
      RECT 768.235 -0.845 768.565 -0.515 ;
      RECT 767.555 -1.525 767.885 -1.195 ;
      RECT 766.875 -0.845 767.205 -0.515 ;
      RECT 766.195 -1.525 766.525 -1.195 ;
      RECT 765.515 -0.845 765.845 -0.515 ;
      RECT 764.835 -1.525 765.165 -1.195 ;
      RECT 764.155 -0.845 764.485 -0.515 ;
      RECT 763.475 -1.525 763.805 -1.195 ;
      RECT 762.795 -0.845 763.125 -0.515 ;
      RECT 762.115 -1.525 762.445 -1.195 ;
      RECT 761.435 -0.845 761.765 -0.515 ;
      RECT 760.755 -1.525 761.085 -1.195 ;
      RECT 760.075 -0.845 760.405 -0.515 ;
      RECT 759.395 -1.525 759.725 -1.195 ;
      RECT 758.715 -0.845 759.045 -0.515 ;
      RECT 758.035 -1.525 758.365 -1.195 ;
      RECT 757.355 -0.845 757.685 -0.515 ;
      RECT 756.675 -1.525 757.005 -1.195 ;
      RECT 755.995 -0.845 756.325 -0.515 ;
      RECT 755.315 -1.525 755.645 -1.195 ;
      RECT 754.635 -0.845 754.965 -0.515 ;
      RECT 753.955 -1.525 754.285 -1.195 ;
      RECT 753.275 -0.845 753.605 -0.515 ;
      RECT 752.595 -1.525 752.925 -1.195 ;
      RECT 751.915 -0.845 752.245 -0.515 ;
      RECT 751.235 -1.525 751.565 -1.195 ;
      RECT 750.555 -0.845 750.885 -0.515 ;
      RECT 749.875 -1.525 750.205 -1.195 ;
      RECT 749.195 -0.845 749.525 -0.515 ;
      RECT 748.515 -1.525 748.845 -1.195 ;
      RECT 747.835 -0.845 748.165 -0.515 ;
      RECT 747.155 -1.525 747.485 -1.195 ;
      RECT 746.475 -0.845 746.805 -0.515 ;
      RECT 745.795 -1.525 746.125 -1.195 ;
      RECT 745.115 -0.845 745.445 -0.515 ;
      RECT 744.435 -1.525 744.765 -1.195 ;
      RECT 743.755 -0.845 744.085 -0.515 ;
      RECT 743.075 -1.525 743.405 -1.195 ;
      RECT 742.395 -0.845 742.725 -0.515 ;
      RECT 741.715 -1.525 742.045 -1.195 ;
      RECT 741.035 -0.845 741.365 -0.515 ;
      RECT 740.355 -1.525 740.685 -1.195 ;
      RECT 739.675 -0.845 740.005 -0.515 ;
      RECT 738.995 -1.525 739.325 -1.195 ;
      RECT 738.315 -0.845 738.645 -0.515 ;
      RECT 737.635 -1.525 737.965 -1.195 ;
      RECT 736.955 -0.845 737.285 -0.515 ;
      RECT 736.275 -1.525 736.605 -1.195 ;
      RECT 735.595 -0.845 735.925 -0.515 ;
      RECT 734.915 -1.525 735.245 -1.195 ;
      RECT 734.235 -0.845 734.565 -0.515 ;
      RECT 733.555 -1.525 733.885 -1.195 ;
      RECT 732.875 -0.845 733.205 -0.515 ;
      RECT 732.195 -1.525 732.525 -1.195 ;
      RECT 731.515 -0.845 731.845 -0.515 ;
      RECT 730.835 -1.525 731.165 -1.195 ;
      RECT 730.155 -0.845 730.485 -0.515 ;
      RECT 729.475 -1.525 729.805 -1.195 ;
      RECT 728.795 -0.845 729.125 -0.515 ;
      RECT 728.115 -1.525 728.445 -1.195 ;
      RECT 727.435 -0.845 727.765 -0.515 ;
      RECT 726.755 -1.525 727.085 -1.195 ;
      RECT 726.075 -0.845 726.405 -0.515 ;
      RECT 725.395 -1.525 725.725 -1.195 ;
      RECT 724.715 -0.845 725.045 -0.515 ;
      RECT 724.035 -1.525 724.365 -1.195 ;
      RECT 723.355 -0.845 723.685 -0.515 ;
      RECT 722.675 -1.525 723.005 -1.195 ;
      RECT 721.995 -0.845 722.325 -0.515 ;
      RECT 721.315 -1.525 721.645 -1.195 ;
      RECT 720.635 -0.845 720.965 -0.515 ;
      RECT 719.955 -1.525 720.285 -1.195 ;
      RECT 719.275 -0.845 719.605 -0.515 ;
      RECT 718.595 -1.525 718.925 -1.195 ;
      RECT 717.915 -0.845 718.245 -0.515 ;
      RECT 717.235 -1.525 717.565 -1.195 ;
      RECT 716.555 -0.845 716.885 -0.515 ;
      RECT 715.875 -1.525 716.205 -1.195 ;
      RECT 715.195 -0.845 715.525 -0.515 ;
      RECT 714.515 -1.525 714.845 -1.195 ;
      RECT 713.835 -0.845 714.165 -0.515 ;
      RECT 713.155 -1.525 713.485 -1.195 ;
      RECT 712.475 -0.845 712.805 -0.515 ;
      RECT 711.795 -1.525 712.125 -1.195 ;
      RECT 711.115 -0.845 711.445 -0.515 ;
      RECT 710.435 -1.525 710.765 -1.195 ;
      RECT 709.755 -0.845 710.085 -0.515 ;
      RECT 709.075 -1.525 709.405 -1.195 ;
      RECT 708.395 -0.845 708.725 -0.515 ;
      RECT 707.715 -1.525 708.045 -1.195 ;
      RECT 707.035 -0.845 707.365 -0.515 ;
      RECT 706.355 -1.525 706.685 -1.195 ;
      RECT 705.675 -0.845 706.005 -0.515 ;
      RECT 704.995 -1.525 705.325 -1.195 ;
      RECT 704.315 -0.845 704.645 -0.515 ;
      RECT 703.635 -1.525 703.965 -1.195 ;
      RECT 702.955 -0.845 703.285 -0.515 ;
      RECT 702.275 -1.525 702.605 -1.195 ;
      RECT 701.595 -0.845 701.925 -0.515 ;
      RECT 700.915 -1.525 701.245 -1.195 ;
      RECT 700.235 -0.845 700.565 -0.515 ;
      RECT 699.555 -1.525 699.885 -1.195 ;
      RECT 698.875 -0.845 699.205 -0.515 ;
      RECT 698.195 -1.525 698.525 -1.195 ;
      RECT 697.515 -0.845 697.845 -0.515 ;
      RECT 696.835 -1.525 697.165 -1.195 ;
      RECT 696.155 -0.845 696.485 -0.515 ;
      RECT 695.475 -1.525 695.805 -1.195 ;
      RECT 694.795 -0.845 695.125 -0.515 ;
      RECT 694.115 -1.525 694.445 -1.195 ;
      RECT 693.435 -0.845 693.765 -0.515 ;
      RECT 692.755 -1.525 693.085 -1.195 ;
      RECT 692.075 -0.845 692.405 -0.515 ;
      RECT 691.395 -1.525 691.725 -1.195 ;
      RECT 690.715 -0.845 691.045 -0.515 ;
      RECT 690.035 -1.525 690.365 -1.195 ;
      RECT 689.355 -0.845 689.685 -0.515 ;
      RECT 688.675 -1.525 689.005 -1.195 ;
      RECT 687.995 -0.845 688.325 -0.515 ;
      RECT 687.315 -1.525 687.645 -1.195 ;
      RECT 686.635 -0.845 686.965 -0.515 ;
      RECT 685.955 -1.525 686.285 -1.195 ;
      RECT 685.275 -0.845 685.605 -0.515 ;
      RECT 684.595 -1.525 684.925 -1.195 ;
      RECT 683.915 -0.845 684.245 -0.515 ;
      RECT 683.235 -1.525 683.565 -1.195 ;
      RECT 682.555 -0.845 682.885 -0.515 ;
      RECT 681.875 -1.525 682.205 -1.195 ;
      RECT 681.195 -0.845 681.525 -0.515 ;
      RECT 680.515 -1.525 680.845 -1.195 ;
      RECT 679.835 -0.845 680.165 -0.515 ;
      RECT 679.155 -1.525 679.485 -1.195 ;
      RECT 678.475 -0.845 678.805 -0.515 ;
      RECT 677.795 -1.525 678.125 -1.195 ;
      RECT 677.115 -0.845 677.445 -0.515 ;
      RECT 676.435 -1.525 676.765 -1.195 ;
      RECT 675.755 -0.845 676.085 -0.515 ;
      RECT 675.075 -1.525 675.405 -1.195 ;
      RECT 674.395 -0.845 674.725 -0.515 ;
      RECT 673.715 -1.525 674.045 -1.195 ;
      RECT 673.035 -0.845 673.365 -0.515 ;
      RECT 672.355 -1.525 672.685 -1.195 ;
      RECT 671.675 -0.845 672.005 -0.515 ;
      RECT 670.995 -1.525 671.325 -1.195 ;
      RECT 670.315 -0.845 670.645 -0.515 ;
      RECT 669.635 -1.525 669.965 -1.195 ;
      RECT 668.955 -0.845 669.285 -0.515 ;
      RECT 668.275 -1.525 668.605 -1.195 ;
      RECT 667.595 -0.845 667.925 -0.515 ;
      RECT 666.915 -1.525 667.245 -1.195 ;
      RECT 666.235 -0.845 666.565 -0.515 ;
      RECT 665.555 -1.525 665.885 -1.195 ;
      RECT 664.875 -0.845 665.205 -0.515 ;
      RECT 664.195 -1.525 664.525 -1.195 ;
      RECT 663.515 -0.845 663.845 -0.515 ;
      RECT 662.835 -1.525 663.165 -1.195 ;
      RECT 662.155 -0.845 662.485 -0.515 ;
      RECT 661.475 -1.525 661.805 -1.195 ;
      RECT 660.795 -0.845 661.125 -0.515 ;
      RECT 660.115 -1.525 660.445 -1.195 ;
      RECT 659.435 -0.845 659.765 -0.515 ;
      RECT 658.755 -1.525 659.085 -1.195 ;
      RECT 658.075 -0.845 658.405 -0.515 ;
      RECT 657.395 -1.525 657.725 -1.195 ;
      RECT 656.715 -0.845 657.045 -0.515 ;
      RECT 656.035 -1.525 656.365 -1.195 ;
      RECT 655.355 -0.845 655.685 -0.515 ;
      RECT 654.675 -1.525 655.005 -1.195 ;
      RECT 653.995 -0.845 654.325 -0.515 ;
      RECT 653.315 -1.525 653.645 -1.195 ;
      RECT 652.635 -0.845 652.965 -0.515 ;
      RECT 651.955 -1.525 652.285 -1.195 ;
      RECT 651.275 -0.845 651.605 -0.515 ;
      RECT 650.595 -1.525 650.925 -1.195 ;
      RECT 649.915 -0.845 650.245 -0.515 ;
      RECT 649.235 -1.525 649.565 -1.195 ;
      RECT 648.555 -0.845 648.885 -0.515 ;
      RECT 647.875 -1.525 648.205 -1.195 ;
      RECT 647.195 -0.845 647.525 -0.515 ;
      RECT 646.515 -1.525 646.845 -1.195 ;
      RECT 645.835 -0.845 646.165 -0.515 ;
      RECT 645.155 -1.525 645.485 -1.195 ;
      RECT 644.475 -0.845 644.805 -0.515 ;
      RECT 643.795 -1.525 644.125 -1.195 ;
      RECT 643.115 -0.845 643.445 -0.515 ;
      RECT 642.435 -1.525 642.765 -1.195 ;
      RECT 641.755 -0.845 642.085 -0.515 ;
      RECT 641.075 -1.525 641.405 -1.195 ;
      RECT 640.395 -0.845 640.725 -0.515 ;
      RECT 639.715 -1.525 640.045 -1.195 ;
      RECT 639.035 -0.845 639.365 -0.515 ;
      RECT 638.355 -1.525 638.685 -1.195 ;
      RECT 637.675 -0.845 638.005 -0.515 ;
      RECT 636.995 -1.525 637.325 -1.195 ;
      RECT 636.315 -0.845 636.645 -0.515 ;
      RECT 635.635 -1.525 635.965 -1.195 ;
      RECT 634.955 -0.845 635.285 -0.515 ;
      RECT 634.275 -1.525 634.605 -1.195 ;
      RECT 633.595 -0.845 633.925 -0.515 ;
      RECT 632.915 -1.525 633.245 -1.195 ;
      RECT 632.235 -0.845 632.565 -0.515 ;
      RECT 631.555 -1.525 631.885 -1.195 ;
      RECT 630.875 -0.845 631.205 -0.515 ;
      RECT 630.195 -1.525 630.525 -1.195 ;
      RECT 629.515 -0.845 629.845 -0.515 ;
      RECT 628.835 -1.525 629.165 -1.195 ;
      RECT 628.155 -0.845 628.485 -0.515 ;
      RECT 627.475 -1.525 627.805 -1.195 ;
      RECT 626.795 -0.845 627.125 -0.515 ;
      RECT 626.115 -1.525 626.445 -1.195 ;
      RECT 625.435 -0.845 625.765 -0.515 ;
      RECT 624.755 -1.525 625.085 -1.195 ;
      RECT 624.075 -0.845 624.405 -0.515 ;
      RECT 623.395 -1.525 623.725 -1.195 ;
      RECT 622.715 -0.845 623.045 -0.515 ;
      RECT 622.035 -1.525 622.365 -1.195 ;
      RECT 621.355 -0.845 621.685 -0.515 ;
      RECT 620.675 -1.525 621.005 -1.195 ;
      RECT 619.995 -0.845 620.325 -0.515 ;
      RECT 619.315 -1.525 619.645 -1.195 ;
      RECT 618.635 -0.845 618.965 -0.515 ;
      RECT 617.955 -1.525 618.285 -1.195 ;
      RECT 617.275 -0.845 617.605 -0.515 ;
      RECT 616.595 -1.525 616.925 -1.195 ;
      RECT 615.915 -0.845 616.245 -0.515 ;
      RECT 615.235 -1.525 615.565 -1.195 ;
      RECT 614.555 -0.845 614.885 -0.515 ;
      RECT 613.875 -1.525 614.205 -1.195 ;
      RECT 613.195 -0.845 613.525 -0.515 ;
      RECT 612.515 -1.525 612.845 -1.195 ;
      RECT 611.835 -0.845 612.165 -0.515 ;
      RECT 611.155 -1.525 611.485 -1.195 ;
      RECT 610.475 -0.845 610.805 -0.515 ;
      RECT 609.795 -1.525 610.125 -1.195 ;
      RECT 609.115 -0.845 609.445 -0.515 ;
      RECT 608.435 -1.525 608.765 -1.195 ;
      RECT 607.755 -0.845 608.085 -0.515 ;
      RECT 607.075 -1.525 607.405 -1.195 ;
      RECT 606.395 -0.845 606.725 -0.515 ;
      RECT 605.715 -1.525 606.045 -1.195 ;
      RECT 605.035 -0.845 605.365 -0.515 ;
      RECT 604.355 -1.525 604.685 -1.195 ;
      RECT 603.675 -0.845 604.005 -0.515 ;
      RECT 602.995 -1.525 603.325 -1.195 ;
      RECT 602.315 -0.845 602.645 -0.515 ;
      RECT 601.635 -1.525 601.965 -1.195 ;
      RECT 600.955 -0.845 601.285 -0.515 ;
      RECT 600.275 -1.525 600.605 -1.195 ;
      RECT 599.595 -0.845 599.925 -0.515 ;
      RECT 598.915 -1.525 599.245 -1.195 ;
      RECT 598.235 -0.845 598.565 -0.515 ;
      RECT 597.555 -1.525 597.885 -1.195 ;
      RECT 596.875 -0.845 597.205 -0.515 ;
      RECT 596.195 -1.525 596.525 -1.195 ;
      RECT 595.515 -0.845 595.845 -0.515 ;
      RECT 594.835 -1.525 595.165 -1.195 ;
      RECT 594.155 -0.845 594.485 -0.515 ;
      RECT 593.475 -1.525 593.805 -1.195 ;
      RECT 592.795 -0.845 593.125 -0.515 ;
      RECT 592.115 -1.525 592.445 -1.195 ;
      RECT 591.435 -0.845 591.765 -0.515 ;
      RECT 590.755 -1.525 591.085 -1.195 ;
      RECT 590.075 -0.845 590.405 -0.515 ;
      RECT 589.395 -1.525 589.725 -1.195 ;
      RECT 588.715 -0.845 589.045 -0.515 ;
      RECT 588.035 -1.525 588.365 -1.195 ;
      RECT 587.355 -0.845 587.685 -0.515 ;
      RECT 586.675 -1.525 587.005 -1.195 ;
      RECT 585.995 -0.845 586.325 -0.515 ;
      RECT 585.315 -1.525 585.645 -1.195 ;
      RECT 584.635 -0.845 584.965 -0.515 ;
      RECT 583.955 -1.525 584.285 -1.195 ;
      RECT 583.275 -0.845 583.605 -0.515 ;
      RECT 582.595 -1.525 582.925 -1.195 ;
      RECT 581.915 -0.845 582.245 -0.515 ;
      RECT 581.235 -1.525 581.565 -1.195 ;
      RECT 580.555 -0.845 580.885 -0.515 ;
      RECT 579.875 -1.525 580.205 -1.195 ;
      RECT 579.195 -0.845 579.525 -0.515 ;
      RECT 578.515 -1.525 578.845 -1.195 ;
      RECT 577.835 -0.845 578.165 -0.515 ;
      RECT 577.155 -1.525 577.485 -1.195 ;
      RECT 576.475 -0.845 576.805 -0.515 ;
      RECT 575.795 -1.525 576.125 -1.195 ;
      RECT 575.115 -0.845 575.445 -0.515 ;
      RECT 574.435 -1.525 574.765 -1.195 ;
      RECT 573.755 -0.845 574.085 -0.515 ;
      RECT 573.075 -1.525 573.405 -1.195 ;
      RECT 572.395 -0.845 572.725 -0.515 ;
      RECT 571.715 -1.525 572.045 -1.195 ;
      RECT 571.035 -0.845 571.365 -0.515 ;
      RECT 570.355 -1.525 570.685 -1.195 ;
      RECT 569.675 -0.845 570.005 -0.515 ;
      RECT 568.995 -1.525 569.325 -1.195 ;
      RECT 568.315 -0.845 568.645 -0.515 ;
      RECT 567.635 -1.525 567.965 -1.195 ;
      RECT 566.955 -0.845 567.285 -0.515 ;
      RECT 566.275 -1.525 566.605 -1.195 ;
      RECT 565.595 -0.845 565.925 -0.515 ;
      RECT 564.915 -1.525 565.245 -1.195 ;
      RECT 564.235 -0.845 564.565 -0.515 ;
      RECT 563.555 -1.525 563.885 -1.195 ;
      RECT 562.875 -0.845 563.205 -0.515 ;
      RECT 562.195 -1.525 562.525 -1.195 ;
      RECT 561.515 -0.845 561.845 -0.515 ;
      RECT 560.835 -1.525 561.165 -1.195 ;
      RECT 560.155 -0.845 560.485 -0.515 ;
      RECT 559.475 -1.525 559.805 -1.195 ;
      RECT 558.795 -0.845 559.125 -0.515 ;
      RECT 558.115 -1.525 558.445 -1.195 ;
      RECT 557.435 -0.845 557.765 -0.515 ;
      RECT 556.755 -1.525 557.085 -1.195 ;
      RECT 556.075 -0.845 556.405 -0.515 ;
      RECT 555.395 -1.525 555.725 -1.195 ;
      RECT 554.715 -0.845 555.045 -0.515 ;
      RECT 554.035 -1.525 554.365 -1.195 ;
      RECT 553.355 -0.845 553.685 -0.515 ;
      RECT 552.675 -1.525 553.005 -1.195 ;
      RECT 551.995 -0.845 552.325 -0.515 ;
      RECT 551.315 -1.525 551.645 -1.195 ;
      RECT 550.635 -0.845 550.965 -0.515 ;
      RECT 549.955 -1.525 550.285 -1.195 ;
      RECT 549.275 -0.845 549.605 -0.515 ;
      RECT 548.595 -1.525 548.925 -1.195 ;
      RECT 547.915 -0.845 548.245 -0.515 ;
      RECT 547.235 -1.525 547.565 -1.195 ;
      RECT 546.555 -0.845 546.885 -0.515 ;
      RECT 545.875 -1.525 546.205 -1.195 ;
      RECT 545.195 -0.845 545.525 -0.515 ;
      RECT 544.515 -1.525 544.845 -1.195 ;
      RECT 543.835 -0.845 544.165 -0.515 ;
      RECT 543.155 -1.525 543.485 -1.195 ;
      RECT 542.475 -0.845 542.805 -0.515 ;
      RECT 541.795 -1.525 542.125 -1.195 ;
      RECT 541.115 -0.845 541.445 -0.515 ;
      RECT 540.435 -1.525 540.765 -1.195 ;
      RECT 539.755 -0.845 540.085 -0.515 ;
      RECT 539.075 -1.525 539.405 -1.195 ;
      RECT 538.395 -0.845 538.725 -0.515 ;
      RECT 537.715 -1.525 538.045 -1.195 ;
      RECT 537.035 -0.845 537.365 -0.515 ;
      RECT 536.355 -1.525 536.685 -1.195 ;
      RECT 535.675 -0.845 536.005 -0.515 ;
      RECT 534.995 -1.525 535.325 -1.195 ;
      RECT 534.315 -0.845 534.645 -0.515 ;
      RECT 533.635 -1.525 533.965 -1.195 ;
      RECT 532.955 -0.845 533.285 -0.515 ;
      RECT 532.275 -1.525 532.605 -1.195 ;
      RECT 531.595 -0.845 531.925 -0.515 ;
      RECT 530.915 -1.525 531.245 -1.195 ;
      RECT 530.235 -0.845 530.565 -0.515 ;
      RECT 529.555 -1.525 529.885 -1.195 ;
      RECT 528.875 -0.845 529.205 -0.515 ;
      RECT 528.195 -1.525 528.525 -1.195 ;
      RECT 527.515 -0.845 527.845 -0.515 ;
      RECT 526.835 -1.525 527.165 -1.195 ;
      RECT 526.155 -0.845 526.485 -0.515 ;
      RECT 525.475 -1.525 525.805 -1.195 ;
      RECT 524.795 -0.845 525.125 -0.515 ;
      RECT 524.115 -1.525 524.445 -1.195 ;
      RECT 523.435 -0.845 523.765 -0.515 ;
      RECT 522.755 -1.525 523.085 -1.195 ;
      RECT 522.075 -0.845 522.405 -0.515 ;
      RECT 521.395 -1.525 521.725 -1.195 ;
      RECT 520.715 -0.845 521.045 -0.515 ;
      RECT 520.035 -1.525 520.365 -1.195 ;
      RECT 519.355 -0.845 519.685 -0.515 ;
      RECT 518.675 -1.525 519.005 -1.195 ;
      RECT 517.995 -0.845 518.325 -0.515 ;
      RECT 517.315 -1.525 517.645 -1.195 ;
      RECT 516.635 -0.845 516.965 -0.515 ;
      RECT 515.955 -1.525 516.285 -1.195 ;
      RECT 515.275 -0.845 515.605 -0.515 ;
      RECT 514.595 -1.525 514.925 -1.195 ;
      RECT 513.915 -0.845 514.245 -0.515 ;
      RECT 513.235 -1.525 513.565 -1.195 ;
      RECT 512.555 -0.845 512.885 -0.515 ;
      RECT 511.875 -1.525 512.205 -1.195 ;
      RECT 511.195 -0.845 511.525 -0.515 ;
      RECT 510.515 -1.525 510.845 -1.195 ;
      RECT 509.835 -0.845 510.165 -0.515 ;
      RECT 509.155 -1.525 509.485 -1.195 ;
      RECT 508.475 -0.845 508.805 -0.515 ;
      RECT 507.795 -1.525 508.125 -1.195 ;
      RECT 507.115 -0.845 507.445 -0.515 ;
      RECT 506.435 -1.525 506.765 -1.195 ;
      RECT 505.755 -0.845 506.085 -0.515 ;
      RECT 505.075 -1.525 505.405 -1.195 ;
      RECT 504.395 -0.845 504.725 -0.515 ;
      RECT 503.715 -1.525 504.045 -1.195 ;
      RECT 503.035 -0.845 503.365 -0.515 ;
      RECT 502.355 -1.525 502.685 -1.195 ;
      RECT 501.675 -0.845 502.005 -0.515 ;
      RECT 500.995 -1.525 501.325 -1.195 ;
      RECT 500.315 -0.845 500.645 -0.515 ;
      RECT 499.635 -1.525 499.965 -1.195 ;
      RECT 498.955 -0.845 499.285 -0.515 ;
      RECT 498.275 -1.525 498.605 -1.195 ;
      RECT 497.595 -0.845 497.925 -0.515 ;
      RECT 496.915 -1.525 497.245 -1.195 ;
      RECT 496.235 -0.845 496.565 -0.515 ;
      RECT 495.555 -1.525 495.885 -1.195 ;
      RECT 494.875 -0.845 495.205 -0.515 ;
      RECT 494.195 -1.525 494.525 -1.195 ;
      RECT 493.515 -0.845 493.845 -0.515 ;
      RECT 492.835 -1.525 493.165 -1.195 ;
      RECT 492.155 -0.845 492.485 -0.515 ;
      RECT 491.475 -1.525 491.805 -1.195 ;
      RECT 490.795 -0.845 491.125 -0.515 ;
      RECT 490.115 -1.525 490.445 -1.195 ;
      RECT 489.435 -0.845 489.765 -0.515 ;
      RECT 488.755 -1.525 489.085 -1.195 ;
      RECT 488.075 -0.845 488.405 -0.515 ;
      RECT 487.395 -1.525 487.725 -1.195 ;
      RECT 486.715 -0.845 487.045 -0.515 ;
      RECT 486.035 -1.525 486.365 -1.195 ;
      RECT 485.355 -0.845 485.685 -0.515 ;
      RECT 484.675 -1.525 485.005 -1.195 ;
      RECT 483.995 -0.845 484.325 -0.515 ;
      RECT 483.315 -1.525 483.645 -1.195 ;
      RECT 482.635 -0.845 482.965 -0.515 ;
      RECT 481.955 -1.525 482.285 -1.195 ;
      RECT 481.275 -0.845 481.605 -0.515 ;
      RECT 480.595 -1.525 480.925 -1.195 ;
      RECT 479.915 -0.845 480.245 -0.515 ;
      RECT 479.235 -1.525 479.565 -1.195 ;
      RECT 478.555 -0.845 478.885 -0.515 ;
      RECT 477.875 -1.525 478.205 -1.195 ;
      RECT 477.195 -0.845 477.525 -0.515 ;
      RECT 476.515 -1.525 476.845 -1.195 ;
      RECT 475.835 -0.845 476.165 -0.515 ;
      RECT 475.155 -1.525 475.485 -1.195 ;
      RECT 474.475 -0.845 474.805 -0.515 ;
      RECT 473.795 -1.525 474.125 -1.195 ;
      RECT 473.115 -0.845 473.445 -0.515 ;
      RECT 472.435 -1.525 472.765 -1.195 ;
      RECT 471.755 -0.845 472.085 -0.515 ;
      RECT 471.075 -1.525 471.405 -1.195 ;
      RECT 470.395 -0.845 470.725 -0.515 ;
      RECT 469.715 -1.525 470.045 -1.195 ;
      RECT 469.035 -0.845 469.365 -0.515 ;
      RECT 468.355 -1.525 468.685 -1.195 ;
      RECT 467.675 -0.845 468.005 -0.515 ;
      RECT 466.995 -1.525 467.325 -1.195 ;
      RECT 466.315 -0.845 466.645 -0.515 ;
      RECT 465.635 -1.525 465.965 -1.195 ;
      RECT 464.955 -0.845 465.285 -0.515 ;
      RECT 464.275 -1.525 464.605 -1.195 ;
      RECT 463.595 -0.845 463.925 -0.515 ;
      RECT 462.915 -1.525 463.245 -1.195 ;
      RECT 462.235 -0.845 462.565 -0.515 ;
      RECT 461.555 -1.525 461.885 -1.195 ;
      RECT 460.875 -0.845 461.205 -0.515 ;
      RECT 460.195 -1.525 460.525 -1.195 ;
      RECT 459.515 -0.845 459.845 -0.515 ;
      RECT 458.835 -1.525 459.165 -1.195 ;
      RECT 458.155 -0.845 458.485 -0.515 ;
      RECT 457.475 -1.525 457.805 -1.195 ;
      RECT 456.795 -0.845 457.125 -0.515 ;
      RECT 456.115 -1.525 456.445 -1.195 ;
      RECT 455.435 -0.845 455.765 -0.515 ;
      RECT 454.755 -1.525 455.085 -1.195 ;
      RECT 454.075 -0.845 454.405 -0.515 ;
      RECT 453.395 -1.525 453.725 -1.195 ;
      RECT 452.715 -0.845 453.045 -0.515 ;
      RECT 452.035 -1.525 452.365 -1.195 ;
      RECT 451.355 -0.845 451.685 -0.515 ;
      RECT 450.675 -1.525 451.005 -1.195 ;
      RECT 449.995 -0.845 450.325 -0.515 ;
      RECT 449.315 -1.525 449.645 -1.195 ;
      RECT 448.635 -0.845 448.965 -0.515 ;
      RECT 447.955 -1.525 448.285 -1.195 ;
      RECT 447.275 -0.845 447.605 -0.515 ;
      RECT 446.595 -1.525 446.925 -1.195 ;
      RECT 445.915 -0.845 446.245 -0.515 ;
      RECT 445.235 -1.525 445.565 -1.195 ;
      RECT 444.555 -0.845 444.885 -0.515 ;
      RECT 443.875 -1.525 444.205 -1.195 ;
      RECT 443.195 -0.845 443.525 -0.515 ;
      RECT 442.515 -1.525 442.845 -1.195 ;
      RECT 441.835 -0.845 442.165 -0.515 ;
      RECT 441.155 -1.525 441.485 -1.195 ;
      RECT 440.475 -0.845 440.805 -0.515 ;
      RECT 439.795 -1.525 440.125 -1.195 ;
      RECT 439.115 -0.845 439.445 -0.515 ;
      RECT 438.435 -1.525 438.765 -1.195 ;
      RECT 437.755 -0.845 438.085 -0.515 ;
      RECT 437.075 -1.525 437.405 -1.195 ;
      RECT 436.395 -0.845 436.725 -0.515 ;
      RECT 435.715 -1.525 436.045 -1.195 ;
      RECT 435.035 -0.845 435.365 -0.515 ;
      RECT 434.355 -1.525 434.685 -1.195 ;
      RECT 433.675 -0.845 434.005 -0.515 ;
      RECT 432.995 -1.525 433.325 -1.195 ;
      RECT 432.315 -0.845 432.645 -0.515 ;
      RECT 431.635 -1.525 431.965 -1.195 ;
      RECT 430.955 -0.845 431.285 -0.515 ;
      RECT 430.275 -1.525 430.605 -1.195 ;
      RECT 429.595 -0.845 429.925 -0.515 ;
      RECT 428.915 -1.525 429.245 -1.195 ;
      RECT 428.235 -0.845 428.565 -0.515 ;
      RECT 427.555 -1.525 427.885 -1.195 ;
      RECT 426.875 -0.845 427.205 -0.515 ;
      RECT 426.195 -1.525 426.525 -1.195 ;
      RECT 425.515 -0.845 425.845 -0.515 ;
      RECT 424.835 -1.525 425.165 -1.195 ;
      RECT 424.155 -0.845 424.485 -0.515 ;
      RECT 423.475 -1.525 423.805 -1.195 ;
      RECT 422.795 -0.845 423.125 -0.515 ;
      RECT 422.115 -1.525 422.445 -1.195 ;
      RECT 421.435 -0.845 421.765 -0.515 ;
      RECT 420.755 -1.525 421.085 -1.195 ;
      RECT 420.075 -0.845 420.405 -0.515 ;
      RECT 419.395 -1.525 419.725 -1.195 ;
      RECT 418.715 -0.845 419.045 -0.515 ;
      RECT 418.035 -1.525 418.365 -1.195 ;
      RECT 417.355 -0.845 417.685 -0.515 ;
      RECT 416.675 -1.525 417.005 -1.195 ;
      RECT 415.995 -0.845 416.325 -0.515 ;
      RECT 415.315 -1.525 415.645 -1.195 ;
      RECT 414.635 -0.845 414.965 -0.515 ;
      RECT 413.955 -1.525 414.285 -1.195 ;
      RECT 413.275 -0.845 413.605 -0.515 ;
      RECT 412.595 -1.525 412.925 -1.195 ;
      RECT 411.915 -0.845 412.245 -0.515 ;
      RECT 411.235 -1.525 411.565 -1.195 ;
      RECT 410.555 -0.845 410.885 -0.515 ;
      RECT 409.875 -1.525 410.205 -1.195 ;
      RECT 409.195 -0.845 409.525 -0.515 ;
      RECT 408.515 -1.525 408.845 -1.195 ;
      RECT 407.835 -0.845 408.165 -0.515 ;
      RECT 407.155 -1.525 407.485 -1.195 ;
      RECT 406.475 -0.845 406.805 -0.515 ;
      RECT 405.795 -1.525 406.125 -1.195 ;
      RECT 405.115 -0.845 405.445 -0.515 ;
      RECT 404.435 -1.525 404.765 -1.195 ;
      RECT 403.755 -0.845 404.085 -0.515 ;
      RECT 403.075 -1.525 403.405 -1.195 ;
      RECT 402.395 -0.845 402.725 -0.515 ;
      RECT 401.715 -1.525 402.045 -1.195 ;
      RECT 401.035 -0.845 401.365 -0.515 ;
      RECT 400.355 -1.525 400.685 -1.195 ;
      RECT 399.675 -0.845 400.005 -0.515 ;
      RECT 398.995 -1.525 399.325 -1.195 ;
      RECT 398.315 -0.845 398.645 -0.515 ;
      RECT 397.635 -1.525 397.965 -1.195 ;
      RECT 396.955 -0.845 397.285 -0.515 ;
      RECT 396.275 -1.525 396.605 -1.195 ;
      RECT 395.595 -0.845 395.925 -0.515 ;
      RECT 394.915 -1.525 395.245 -1.195 ;
      RECT 394.235 -0.845 394.565 -0.515 ;
      RECT 393.555 -1.525 393.885 -1.195 ;
      RECT 392.875 -0.845 393.205 -0.515 ;
      RECT 392.195 -1.525 392.525 -1.195 ;
      RECT 391.515 -0.845 391.845 -0.515 ;
      RECT 390.835 -1.525 391.165 -1.195 ;
      RECT 390.155 -0.845 390.485 -0.515 ;
      RECT 389.475 -1.525 389.805 -1.195 ;
      RECT 388.795 -0.845 389.125 -0.515 ;
      RECT 388.115 -1.525 388.445 -1.195 ;
      RECT 387.435 -0.845 387.765 -0.515 ;
      RECT 386.755 -1.525 387.085 -1.195 ;
      RECT 386.075 -0.845 386.405 -0.515 ;
      RECT 385.395 -1.525 385.725 -1.195 ;
      RECT 384.715 -0.845 385.045 -0.515 ;
      RECT 384.035 -1.525 384.365 -1.195 ;
      RECT 383.355 -0.845 383.685 -0.515 ;
      RECT 382.675 -1.525 383.005 -1.195 ;
      RECT 381.995 -0.845 382.325 -0.515 ;
      RECT 381.315 -1.525 381.645 -1.195 ;
      RECT 380.635 -0.845 380.965 -0.515 ;
      RECT 379.955 -1.525 380.285 -1.195 ;
      RECT 379.275 -0.845 379.605 -0.515 ;
      RECT 378.595 -1.525 378.925 -1.195 ;
      RECT 377.915 -0.845 378.245 -0.515 ;
      RECT 377.235 -1.525 377.565 -1.195 ;
      RECT 376.555 -0.845 376.885 -0.515 ;
      RECT 375.875 -1.525 376.205 -1.195 ;
      RECT 375.195 -0.845 375.525 -0.515 ;
      RECT 374.515 -1.525 374.845 -1.195 ;
      RECT 373.835 -0.845 374.165 -0.515 ;
      RECT 373.155 -1.525 373.485 -1.195 ;
      RECT 372.475 -0.845 372.805 -0.515 ;
      RECT 371.795 -1.525 372.125 -1.195 ;
      RECT 371.115 -0.845 371.445 -0.515 ;
      RECT 370.435 -1.525 370.765 -1.195 ;
      RECT 369.755 -0.845 370.085 -0.515 ;
      RECT 369.075 -1.525 369.405 -1.195 ;
      RECT 368.395 -0.845 368.725 -0.515 ;
      RECT 367.715 -1.525 368.045 -1.195 ;
      RECT 367.035 -0.845 367.365 -0.515 ;
      RECT 366.355 -1.525 366.685 -1.195 ;
      RECT 365.675 -0.845 366.005 -0.515 ;
      RECT 364.995 -1.525 365.325 -1.195 ;
      RECT 364.315 -0.845 364.645 -0.515 ;
      RECT 363.635 -1.525 363.965 -1.195 ;
      RECT 362.955 -0.845 363.285 -0.515 ;
      RECT 362.275 -1.525 362.605 -1.195 ;
      RECT 361.595 -0.845 361.925 -0.515 ;
      RECT 360.915 -1.525 361.245 -1.195 ;
      RECT 360.235 -0.845 360.565 -0.515 ;
      RECT 359.555 -1.525 359.885 -1.195 ;
      RECT 358.875 -0.845 359.205 -0.515 ;
      RECT 358.195 -1.525 358.525 -1.195 ;
      RECT 357.515 -0.845 357.845 -0.515 ;
      RECT 356.835 -1.525 357.165 -1.195 ;
      RECT 356.155 -0.845 356.485 -0.515 ;
      RECT 355.475 -1.525 355.805 -1.195 ;
      RECT 354.795 -0.845 355.125 -0.515 ;
      RECT 354.115 -1.525 354.445 -1.195 ;
      RECT 353.435 -0.845 353.765 -0.515 ;
      RECT 352.755 -1.525 353.085 -1.195 ;
      RECT 352.075 -0.845 352.405 -0.515 ;
      RECT 351.395 -1.525 351.725 -1.195 ;
      RECT 350.715 -0.845 351.045 -0.515 ;
      RECT 350.035 -1.525 350.365 -1.195 ;
      RECT 349.355 -0.845 349.685 -0.515 ;
      RECT 348.675 -1.525 349.005 -1.195 ;
      RECT 347.995 -0.845 348.325 -0.515 ;
      RECT 347.315 -1.525 347.645 -1.195 ;
      RECT 346.635 -0.845 346.965 -0.515 ;
      RECT 345.955 -1.525 346.285 -1.195 ;
      RECT 345.275 -0.845 345.605 -0.515 ;
      RECT 344.595 -1.525 344.925 -1.195 ;
      RECT 343.915 -0.845 344.245 -0.515 ;
      RECT 343.235 -1.525 343.565 -1.195 ;
      RECT 342.555 -0.845 342.885 -0.515 ;
      RECT 341.875 -1.525 342.205 -1.195 ;
      RECT 341.195 -0.845 341.525 -0.515 ;
      RECT 340.515 -1.525 340.845 -1.195 ;
      RECT 339.835 -0.845 340.165 -0.515 ;
      RECT 339.155 -1.525 339.485 -1.195 ;
      RECT 338.475 -0.845 338.805 -0.515 ;
      RECT 337.795 -1.525 338.125 -1.195 ;
      RECT 337.115 -0.845 337.445 -0.515 ;
      RECT 336.435 -1.525 336.765 -1.195 ;
      RECT 335.755 -0.845 336.085 -0.515 ;
      RECT 335.075 -1.525 335.405 -1.195 ;
      RECT 334.395 -0.845 334.725 -0.515 ;
      RECT 333.715 -1.525 334.045 -1.195 ;
      RECT 333.035 -0.845 333.365 -0.515 ;
      RECT 332.355 -1.525 332.685 -1.195 ;
      RECT 331.675 -0.845 332.005 -0.515 ;
      RECT 330.995 -1.525 331.325 -1.195 ;
      RECT 330.315 -0.845 330.645 -0.515 ;
      RECT 329.635 -1.525 329.965 -1.195 ;
      RECT 328.955 -0.845 329.285 -0.515 ;
      RECT 328.275 -1.525 328.605 -1.195 ;
      RECT 327.595 -0.845 327.925 -0.515 ;
      RECT 326.915 -1.525 327.245 -1.195 ;
      RECT 326.235 -0.845 326.565 -0.515 ;
      RECT 325.555 -1.525 325.885 -1.195 ;
      RECT 324.875 -0.845 325.205 -0.515 ;
      RECT 324.195 -1.525 324.525 -1.195 ;
      RECT 323.515 -0.845 323.845 -0.515 ;
      RECT 322.835 -1.525 323.165 -1.195 ;
      RECT 322.155 -0.845 322.485 -0.515 ;
      RECT 321.475 -1.525 321.805 -1.195 ;
      RECT 320.795 -0.845 321.125 -0.515 ;
      RECT 320.115 -1.525 320.445 -1.195 ;
      RECT 319.435 -0.845 319.765 -0.515 ;
      RECT 318.755 -1.525 319.085 -1.195 ;
      RECT 318.075 -0.845 318.405 -0.515 ;
      RECT 317.395 -1.525 317.725 -1.195 ;
      RECT 316.715 -0.845 317.045 -0.515 ;
      RECT 316.035 -1.525 316.365 -1.195 ;
      RECT 315.355 -0.845 315.685 -0.515 ;
      RECT 314.675 -1.525 315.005 -1.195 ;
      RECT 313.995 -0.845 314.325 -0.515 ;
      RECT 313.315 -1.525 313.645 -1.195 ;
      RECT 312.635 -0.845 312.965 -0.515 ;
      RECT 311.955 -1.525 312.285 -1.195 ;
      RECT 311.275 -0.845 311.605 -0.515 ;
      RECT 310.595 -1.525 310.925 -1.195 ;
      RECT 309.915 -0.845 310.245 -0.515 ;
      RECT 309.235 -1.525 309.565 -1.195 ;
      RECT 308.555 -0.845 308.885 -0.515 ;
      RECT 307.875 -1.525 308.205 -1.195 ;
      RECT 307.195 -0.845 307.525 -0.515 ;
      RECT 306.515 -1.525 306.845 -1.195 ;
      RECT 305.835 -0.845 306.165 -0.515 ;
      RECT 305.155 -1.525 305.485 -1.195 ;
      RECT 304.475 -0.845 304.805 -0.515 ;
      RECT 303.795 -1.525 304.125 -1.195 ;
      RECT 303.115 -0.845 303.445 -0.515 ;
      RECT 302.435 -1.525 302.765 -1.195 ;
      RECT 301.755 -0.845 302.085 -0.515 ;
      RECT 301.075 -1.525 301.405 -1.195 ;
      RECT 300.395 -0.845 300.725 -0.515 ;
      RECT 299.715 -1.525 300.045 -1.195 ;
      RECT 299.035 -0.845 299.365 -0.515 ;
      RECT 298.355 -1.525 298.685 -1.195 ;
      RECT 297.675 -0.845 298.005 -0.515 ;
      RECT 296.995 -1.525 297.325 -1.195 ;
      RECT 296.315 -0.845 296.645 -0.515 ;
      RECT 295.635 -1.525 295.965 -1.195 ;
      RECT 294.955 -0.845 295.285 -0.515 ;
      RECT 294.275 -1.525 294.605 -1.195 ;
      RECT 293.595 -0.845 293.925 -0.515 ;
      RECT 292.915 -1.525 293.245 -1.195 ;
      RECT 292.235 -0.845 292.565 -0.515 ;
      RECT 291.555 -1.525 291.885 -1.195 ;
      RECT 290.875 -0.845 291.205 -0.515 ;
      RECT 290.195 -1.525 290.525 -1.195 ;
      RECT 289.515 -0.845 289.845 -0.515 ;
      RECT 288.835 -1.525 289.165 -1.195 ;
      RECT 288.155 -0.845 288.485 -0.515 ;
      RECT 287.475 -1.525 287.805 -1.195 ;
      RECT 286.795 -0.845 287.125 -0.515 ;
      RECT 286.115 -1.525 286.445 -1.195 ;
      RECT 285.435 -0.845 285.765 -0.515 ;
      RECT 284.755 -1.525 285.085 -1.195 ;
      RECT 284.075 -0.845 284.405 -0.515 ;
      RECT 283.395 -1.525 283.725 -1.195 ;
      RECT 282.715 -0.845 283.045 -0.515 ;
      RECT 282.035 -1.525 282.365 -1.195 ;
      RECT 281.355 -0.845 281.685 -0.515 ;
      RECT 280.675 -1.525 281.005 -1.195 ;
      RECT 279.995 -0.845 280.325 -0.515 ;
      RECT 279.315 -1.525 279.645 -1.195 ;
      RECT 278.635 -0.845 278.965 -0.515 ;
      RECT 277.955 -1.525 278.285 -1.195 ;
      RECT 277.275 -0.845 277.605 -0.515 ;
      RECT 276.595 -1.525 276.925 -1.195 ;
      RECT 275.915 -0.845 276.245 -0.515 ;
      RECT 275.235 -1.525 275.565 -1.195 ;
      RECT 274.555 -0.845 274.885 -0.515 ;
      RECT 273.875 -1.525 274.205 -1.195 ;
      RECT 273.195 -0.845 273.525 -0.515 ;
      RECT 272.515 -1.525 272.845 -1.195 ;
      RECT 271.835 -0.845 272.165 -0.515 ;
      RECT 271.155 -1.525 271.485 -1.195 ;
      RECT 270.475 -0.845 270.805 -0.515 ;
      RECT 269.795 -1.525 270.125 -1.195 ;
      RECT 269.115 -0.845 269.445 -0.515 ;
      RECT 268.435 -1.525 268.765 -1.195 ;
      RECT 267.755 -0.845 268.085 -0.515 ;
      RECT 267.075 -1.525 267.405 -1.195 ;
      RECT 266.395 -0.845 266.725 -0.515 ;
      RECT 265.715 -1.525 266.045 -1.195 ;
      RECT 265.035 -0.845 265.365 -0.515 ;
      RECT 264.355 -1.525 264.685 -1.195 ;
      RECT 263.675 -0.845 264.005 -0.515 ;
      RECT 262.995 -1.525 263.325 -1.195 ;
      RECT 262.315 -0.845 262.645 -0.515 ;
      RECT 261.635 -1.525 261.965 -1.195 ;
      RECT 260.955 -0.845 261.285 -0.515 ;
      RECT 260.275 -1.525 260.605 -1.195 ;
      RECT 259.595 -0.845 259.925 -0.515 ;
      RECT 258.915 -1.525 259.245 -1.195 ;
      RECT 258.235 -0.845 258.565 -0.515 ;
      RECT 257.555 -1.525 257.885 -1.195 ;
      RECT 256.875 -0.845 257.205 -0.515 ;
      RECT 256.195 -1.525 256.525 -1.195 ;
      RECT 255.515 -0.845 255.845 -0.515 ;
      RECT 254.835 -1.525 255.165 -1.195 ;
      RECT 254.155 -0.845 254.485 -0.515 ;
      RECT 253.475 -1.525 253.805 -1.195 ;
      RECT 252.795 -0.845 253.125 -0.515 ;
      RECT 252.115 -1.525 252.445 -1.195 ;
      RECT 251.435 -0.845 251.765 -0.515 ;
      RECT 250.755 -1.525 251.085 -1.195 ;
      RECT 250.075 -0.845 250.405 -0.515 ;
      RECT 249.395 -1.525 249.725 -1.195 ;
      RECT 248.715 -0.845 249.045 -0.515 ;
      RECT 248.035 -1.525 248.365 -1.195 ;
      RECT 247.355 -0.845 247.685 -0.515 ;
      RECT 246.675 -1.525 247.005 -1.195 ;
      RECT 245.995 -0.845 246.325 -0.515 ;
      RECT 245.315 -1.525 245.645 -1.195 ;
      RECT 244.635 -0.845 244.965 -0.515 ;
      RECT 243.955 -1.525 244.285 -1.195 ;
      RECT 243.275 -0.845 243.605 -0.515 ;
      RECT 242.595 -1.525 242.925 -1.195 ;
      RECT 241.915 -0.845 242.245 -0.515 ;
      RECT 241.235 -1.525 241.565 -1.195 ;
      RECT 240.555 -0.845 240.885 -0.515 ;
      RECT 239.875 -1.525 240.205 -1.195 ;
      RECT 239.195 -0.845 239.525 -0.515 ;
      RECT 238.515 -1.525 238.845 -1.195 ;
      RECT 237.835 -0.845 238.165 -0.515 ;
      RECT 237.155 -1.525 237.485 -1.195 ;
      RECT 236.475 -0.845 236.805 -0.515 ;
      RECT 235.795 -1.525 236.125 -1.195 ;
      RECT 235.115 -0.845 235.445 -0.515 ;
      RECT 234.435 -1.525 234.765 -1.195 ;
      RECT 233.755 -0.845 234.085 -0.515 ;
      RECT 233.075 -1.525 233.405 -1.195 ;
      RECT 232.395 -0.845 232.725 -0.515 ;
      RECT 231.715 -1.525 232.045 -1.195 ;
      RECT 231.035 -0.845 231.365 -0.515 ;
      RECT 230.355 -1.525 230.685 -1.195 ;
      RECT 229.675 -0.845 230.005 -0.515 ;
      RECT 228.995 -1.525 229.325 -1.195 ;
      RECT 228.315 -0.845 228.645 -0.515 ;
      RECT 227.635 -1.525 227.965 -1.195 ;
      RECT 226.955 -0.845 227.285 -0.515 ;
      RECT 226.275 -1.525 226.605 -1.195 ;
      RECT 225.595 -0.845 225.925 -0.515 ;
      RECT 224.915 -1.525 225.245 -1.195 ;
      RECT 224.235 -0.845 224.565 -0.515 ;
      RECT 223.555 -1.525 223.885 -1.195 ;
      RECT 222.875 -0.845 223.205 -0.515 ;
      RECT 222.195 -1.525 222.525 -1.195 ;
      RECT 221.515 -0.845 221.845 -0.515 ;
      RECT 220.835 -1.525 221.165 -1.195 ;
      RECT 220.155 -0.845 220.485 -0.515 ;
      RECT 219.475 -1.525 219.805 -1.195 ;
      RECT 218.795 -0.845 219.125 -0.515 ;
      RECT 218.115 -1.525 218.445 -1.195 ;
      RECT 217.435 -0.845 217.765 -0.515 ;
      RECT 216.755 -1.525 217.085 -1.195 ;
      RECT 216.075 -0.845 216.405 -0.515 ;
      RECT 215.395 -1.525 215.725 -1.195 ;
      RECT 214.715 -0.845 215.045 -0.515 ;
      RECT 214.035 -1.525 214.365 -1.195 ;
      RECT 213.355 -0.845 213.685 -0.515 ;
      RECT 212.675 -1.525 213.005 -1.195 ;
      RECT 211.995 -0.845 212.325 -0.515 ;
      RECT 211.315 -1.525 211.645 -1.195 ;
      RECT 210.635 -0.845 210.965 -0.515 ;
      RECT 209.955 -1.525 210.285 -1.195 ;
      RECT 209.275 -0.845 209.605 -0.515 ;
      RECT 208.595 -1.525 208.925 -1.195 ;
      RECT 207.915 -0.845 208.245 -0.515 ;
      RECT 207.235 -1.525 207.565 -1.195 ;
      RECT 206.555 -0.845 206.885 -0.515 ;
      RECT 205.875 -1.525 206.205 -1.195 ;
      RECT 205.195 -0.845 205.525 -0.515 ;
      RECT 204.515 -1.525 204.845 -1.195 ;
      RECT 203.835 -0.845 204.165 -0.515 ;
      RECT 203.155 -1.525 203.485 -1.195 ;
      RECT 202.475 -0.845 202.805 -0.515 ;
      RECT 201.795 -1.525 202.125 -1.195 ;
      RECT 201.115 -0.845 201.445 -0.515 ;
      RECT 200.435 -1.525 200.765 -1.195 ;
      RECT 199.755 -0.845 200.085 -0.515 ;
      RECT 199.075 -1.525 199.405 -1.195 ;
      RECT 198.395 -0.845 198.725 -0.515 ;
      RECT 197.715 -1.525 198.045 -1.195 ;
      RECT 197.035 -0.845 197.365 -0.515 ;
      RECT 196.355 -1.525 196.685 -1.195 ;
      RECT 195.675 -0.845 196.005 -0.515 ;
      RECT 194.995 -1.525 195.325 -1.195 ;
      RECT 194.315 -0.845 194.645 -0.515 ;
      RECT 193.635 -1.525 193.965 -1.195 ;
      RECT 192.955 -0.845 193.285 -0.515 ;
      RECT 192.275 -1.525 192.605 -1.195 ;
      RECT 191.595 -0.845 191.925 -0.515 ;
      RECT 190.915 -1.525 191.245 -1.195 ;
      RECT 190.235 -0.845 190.565 -0.515 ;
      RECT 189.555 -1.525 189.885 -1.195 ;
      RECT 188.875 -0.845 189.205 -0.515 ;
      RECT 188.195 -1.525 188.525 -1.195 ;
      RECT 187.515 -0.845 187.845 -0.515 ;
      RECT 186.835 -1.525 187.165 -1.195 ;
      RECT 186.155 -0.845 186.485 -0.515 ;
      RECT 185.475 -1.525 185.805 -1.195 ;
      RECT 184.795 -0.845 185.125 -0.515 ;
      RECT 184.115 -1.525 184.445 -1.195 ;
      RECT 183.435 -0.845 183.765 -0.515 ;
      RECT 182.755 -1.525 183.085 -1.195 ;
      RECT 182.075 -0.845 182.405 -0.515 ;
      RECT 181.395 -1.525 181.725 -1.195 ;
      RECT 180.715 -0.845 181.045 -0.515 ;
      RECT 180.035 -1.525 180.365 -1.195 ;
      RECT 179.355 -0.845 179.685 -0.515 ;
      RECT 178.675 -1.525 179.005 -1.195 ;
      RECT 177.995 -0.845 178.325 -0.515 ;
      RECT 177.315 -1.525 177.645 -1.195 ;
      RECT 176.635 -0.845 176.965 -0.515 ;
      RECT 175.955 -1.525 176.285 -1.195 ;
      RECT 175.275 -0.845 175.605 -0.515 ;
      RECT 174.595 -1.525 174.925 -1.195 ;
      RECT 173.915 -0.845 174.245 -0.515 ;
      RECT 173.235 -1.525 173.565 -1.195 ;
      RECT 172.555 -0.845 172.885 -0.515 ;
      RECT 171.875 -1.525 172.205 -1.195 ;
      RECT 171.195 -0.845 171.525 -0.515 ;
      RECT 170.515 -1.525 170.845 -1.195 ;
      RECT 169.835 -0.845 170.165 -0.515 ;
      RECT 169.155 -1.525 169.485 -1.195 ;
      RECT 168.475 -0.845 168.805 -0.515 ;
      RECT 167.795 -1.525 168.125 -1.195 ;
      RECT 167.115 -0.845 167.445 -0.515 ;
      RECT 166.435 -1.525 166.765 -1.195 ;
      RECT 165.755 -0.845 166.085 -0.515 ;
      RECT 165.075 -1.525 165.405 -1.195 ;
      RECT 164.395 -0.845 164.725 -0.515 ;
      RECT 163.715 -1.525 164.045 -1.195 ;
      RECT 163.035 -0.845 163.365 -0.515 ;
      RECT 162.355 -1.525 162.685 -1.195 ;
      RECT 161.675 -0.845 162.005 -0.515 ;
      RECT 160.995 -1.525 161.325 -1.195 ;
      RECT 160.315 -0.845 160.645 -0.515 ;
      RECT 159.635 -1.525 159.965 -1.195 ;
      RECT 158.955 -0.845 159.285 -0.515 ;
      RECT 158.275 -1.525 158.605 -1.195 ;
      RECT 157.595 -0.845 157.925 -0.515 ;
      RECT 156.915 -1.525 157.245 -1.195 ;
      RECT 156.235 -0.845 156.565 -0.515 ;
      RECT 155.555 -1.525 155.885 -1.195 ;
      RECT 154.875 -0.845 155.205 -0.515 ;
      RECT 154.195 -1.525 154.525 -1.195 ;
      RECT 153.515 -0.845 153.845 -0.515 ;
      RECT 152.835 -1.525 153.165 -1.195 ;
      RECT 152.155 -0.845 152.485 -0.515 ;
      RECT 151.475 -1.525 151.805 -1.195 ;
      RECT 150.795 -0.845 151.125 -0.515 ;
      RECT 150.115 -1.525 150.445 -1.195 ;
      RECT 149.435 -0.845 149.765 -0.515 ;
      RECT 148.755 -1.525 149.085 -1.195 ;
      RECT 148.075 -0.845 148.405 -0.515 ;
      RECT 147.395 -1.525 147.725 -1.195 ;
      RECT 146.715 -0.845 147.045 -0.515 ;
      RECT 146.035 -1.525 146.365 -1.195 ;
      RECT 145.355 -0.845 145.685 -0.515 ;
      RECT 144.675 -1.525 145.005 -1.195 ;
      RECT 143.995 -0.845 144.325 -0.515 ;
      RECT 143.315 -1.525 143.645 -1.195 ;
      RECT 142.635 -0.845 142.965 -0.515 ;
      RECT 141.955 -1.525 142.285 -1.195 ;
      RECT 141.275 -0.845 141.605 -0.515 ;
      RECT 140.595 -1.525 140.925 -1.195 ;
      RECT 139.915 -0.845 140.245 -0.515 ;
      RECT 139.235 -1.525 139.565 -1.195 ;
      RECT 138.555 -0.845 138.885 -0.515 ;
      RECT 137.875 -1.525 138.205 -1.195 ;
      RECT 137.195 -0.845 137.525 -0.515 ;
      RECT 136.515 -1.525 136.845 -1.195 ;
      RECT 135.835 -0.845 136.165 -0.515 ;
      RECT 135.155 -1.525 135.485 -1.195 ;
      RECT 134.475 -0.845 134.805 -0.515 ;
      RECT 133.795 -1.525 134.125 -1.195 ;
      RECT 133.115 -0.845 133.445 -0.515 ;
      RECT 132.435 -1.525 132.765 -1.195 ;
      RECT 131.755 -0.845 132.085 -0.515 ;
      RECT 131.075 -1.525 131.405 -1.195 ;
      RECT 130.395 -0.845 130.725 -0.515 ;
      RECT 129.715 -1.525 130.045 -1.195 ;
      RECT 129.035 -0.845 129.365 -0.515 ;
      RECT 128.355 -1.525 128.685 -1.195 ;
      RECT 127.675 -0.845 128.005 -0.515 ;
      RECT 126.995 -1.525 127.325 -1.195 ;
      RECT 126.315 -0.845 126.645 -0.515 ;
      RECT 125.635 -1.525 125.965 -1.195 ;
      RECT 124.955 -0.845 125.285 -0.515 ;
      RECT 124.275 -1.525 124.605 -1.195 ;
      RECT 123.595 -0.845 123.925 -0.515 ;
      RECT 122.915 -1.525 123.245 -1.195 ;
      RECT 122.235 -0.845 122.565 -0.515 ;
      RECT 121.555 -1.525 121.885 -1.195 ;
      RECT 120.875 -0.845 121.205 -0.515 ;
      RECT 120.195 -1.525 120.525 -1.195 ;
      RECT 119.515 -0.845 119.845 -0.515 ;
      RECT 118.835 -1.525 119.165 -1.195 ;
      RECT 118.155 -0.845 118.485 -0.515 ;
      RECT 117.475 -1.525 117.805 -1.195 ;
      RECT 116.795 -0.845 117.125 -0.515 ;
      RECT 116.115 -1.525 116.445 -1.195 ;
      RECT 115.435 -0.845 115.765 -0.515 ;
      RECT 114.755 -1.525 115.085 -1.195 ;
      RECT 114.075 -0.845 114.405 -0.515 ;
      RECT 113.395 -1.525 113.725 -1.195 ;
      RECT 112.715 -0.845 113.045 -0.515 ;
      RECT 112.035 -1.525 112.365 -1.195 ;
      RECT 111.355 -0.845 111.685 -0.515 ;
      RECT 110.675 -1.525 111.005 -1.195 ;
      RECT 109.995 -0.845 110.325 -0.515 ;
      RECT 109.315 -1.525 109.645 -1.195 ;
      RECT 108.635 -0.845 108.965 -0.515 ;
      RECT 107.955 -1.525 108.285 -1.195 ;
      RECT 107.275 -0.845 107.605 -0.515 ;
      RECT 106.595 -1.525 106.925 -1.195 ;
      RECT 105.915 -0.845 106.245 -0.515 ;
      RECT 105.235 -1.525 105.565 -1.195 ;
      RECT 104.555 -0.845 104.885 -0.515 ;
      RECT 103.875 -1.525 104.205 -1.195 ;
      RECT 103.195 -0.845 103.525 -0.515 ;
      RECT 102.515 -1.525 102.845 -1.195 ;
      RECT 101.835 -0.845 102.165 -0.515 ;
      RECT 101.155 -1.525 101.485 -1.195 ;
      RECT 100.475 -0.845 100.805 -0.515 ;
      RECT 99.795 -1.525 100.125 -1.195 ;
      RECT 99.115 -0.845 99.445 -0.515 ;
      RECT 98.435 -1.525 98.765 -1.195 ;
      RECT 97.755 -0.845 98.085 -0.515 ;
      RECT 97.075 -1.525 97.405 -1.195 ;
      RECT 96.395 -0.845 96.725 -0.515 ;
      RECT 95.715 -1.525 96.045 -1.195 ;
      RECT 95.035 -0.845 95.365 -0.515 ;
      RECT 94.355 -1.525 94.685 -1.195 ;
      RECT 93.675 -0.845 94.005 -0.515 ;
      RECT 92.995 -1.525 93.325 -1.195 ;
      RECT 92.315 -0.845 92.645 -0.515 ;
      RECT 91.635 -1.525 91.965 -1.195 ;
      RECT 90.955 -0.845 91.285 -0.515 ;
      RECT 90.275 -1.525 90.605 -1.195 ;
      RECT 89.595 -0.845 89.925 -0.515 ;
      RECT 88.915 -1.525 89.245 -1.195 ;
      RECT 88.235 -0.845 88.565 -0.515 ;
      RECT 87.555 -1.525 87.885 -1.195 ;
      RECT 86.875 -0.845 87.205 -0.515 ;
      RECT 86.195 -1.525 86.525 -1.195 ;
      RECT 85.515 -0.845 85.845 -0.515 ;
      RECT 84.835 -1.525 85.165 -1.195 ;
      RECT 84.155 -0.845 84.485 -0.515 ;
      RECT 83.475 -1.525 83.805 -1.195 ;
      RECT 82.795 -0.845 83.125 -0.515 ;
      RECT 82.115 -1.525 82.445 -1.195 ;
      RECT 81.435 -0.845 81.765 -0.515 ;
      RECT 80.755 -1.525 81.085 -1.195 ;
      RECT 80.075 -0.845 80.405 -0.515 ;
      RECT 79.395 -1.525 79.725 -1.195 ;
      RECT 78.715 -0.845 79.045 -0.515 ;
      RECT 78.035 -1.525 78.365 -1.195 ;
      RECT 77.355 -0.845 77.685 -0.515 ;
      RECT 76.675 -1.525 77.005 -1.195 ;
      RECT 75.995 -0.845 76.325 -0.515 ;
      RECT 75.315 -1.525 75.645 -1.195 ;
      RECT 74.635 -0.845 74.965 -0.515 ;
      RECT 73.955 -1.525 74.285 -1.195 ;
      RECT 73.275 -0.845 73.605 -0.515 ;
      RECT 72.595 -1.525 72.925 -1.195 ;
      RECT 71.915 -0.845 72.245 -0.515 ;
      RECT 71.235 -1.525 71.565 -1.195 ;
      RECT 70.555 -0.845 70.885 -0.515 ;
      RECT 69.875 -1.525 70.205 -1.195 ;
      RECT 69.195 -0.845 69.525 -0.515 ;
      RECT 68.515 -1.525 68.845 -1.195 ;
      RECT 67.835 -0.845 68.165 -0.515 ;
      RECT 67.155 -1.525 67.485 -1.195 ;
      RECT 66.475 -0.845 66.805 -0.515 ;
      RECT 65.795 -1.525 66.125 -1.195 ;
      RECT 65.115 -0.845 65.445 -0.515 ;
      RECT 64.435 -1.525 64.765 -1.195 ;
      RECT 63.755 -0.845 64.085 -0.515 ;
      RECT 63.075 -1.525 63.405 -1.195 ;
      RECT 62.395 -0.845 62.725 -0.515 ;
      RECT 61.715 -1.525 62.045 -1.195 ;
      RECT 61.035 -0.845 61.365 -0.515 ;
      RECT 60.355 -1.525 60.685 -1.195 ;
      RECT 59.675 -0.845 60.005 -0.515 ;
      RECT 58.995 -1.525 59.325 -1.195 ;
      RECT 58.315 -0.845 58.645 -0.515 ;
      RECT 57.635 -1.525 57.965 -1.195 ;
      RECT 56.955 -0.845 57.285 -0.515 ;
      RECT 56.275 -1.525 56.605 -1.195 ;
      RECT 55.595 -0.845 55.925 -0.515 ;
      RECT 54.915 -1.525 55.245 -1.195 ;
      RECT 54.235 -0.845 54.565 -0.515 ;
      RECT 53.555 -1.525 53.885 -1.195 ;
      RECT 52.875 -0.845 53.205 -0.515 ;
      RECT 52.195 -1.525 52.525 -1.195 ;
      RECT 51.515 -0.845 51.845 -0.515 ;
      RECT 50.835 -1.525 51.165 -1.195 ;
      RECT 50.155 -0.845 50.485 -0.515 ;
      RECT 49.475 -1.525 49.805 -1.195 ;
      RECT 48.795 -0.845 49.125 -0.515 ;
      RECT 48.115 -1.525 48.445 -1.195 ;
      RECT 47.435 -0.845 47.765 -0.515 ;
      RECT 46.755 -1.525 47.085 -1.195 ;
      RECT 46.075 -0.845 46.405 -0.515 ;
      RECT 45.395 -1.525 45.725 -1.195 ;
      RECT 44.715 -0.845 45.045 -0.515 ;
      RECT 44.035 -1.525 44.365 -1.195 ;
      RECT 43.355 -0.845 43.685 -0.515 ;
      RECT 42.675 -1.525 43.005 -1.195 ;
      RECT 41.995 -0.845 42.325 -0.515 ;
      RECT 41.315 -1.525 41.645 -1.195 ;
      RECT 40.635 -0.845 40.965 -0.515 ;
      RECT 39.955 -1.525 40.285 -1.195 ;
      RECT 39.275 -0.845 39.605 -0.515 ;
      RECT 38.595 -1.525 38.925 -1.195 ;
      RECT 37.915 -0.845 38.245 -0.515 ;
      RECT 37.235 -1.525 37.565 -1.195 ;
      RECT 36.555 -0.845 36.885 -0.515 ;
      RECT 35.875 -1.525 36.205 -1.195 ;
      RECT 35.195 -0.845 35.525 -0.515 ;
      RECT 34.515 -1.525 34.845 -1.195 ;
      RECT 33.835 -0.845 34.165 -0.515 ;
      RECT 33.155 -1.525 33.485 -1.195 ;
      RECT 32.475 -0.845 32.805 -0.515 ;
      RECT 31.795 -1.525 32.125 -1.195 ;
      RECT 31.115 -0.845 31.445 -0.515 ;
      RECT 30.435 -1.525 30.765 -1.195 ;
      RECT 29.755 -0.845 30.085 -0.515 ;
      RECT 29.075 -1.525 29.405 -1.195 ;
      RECT 28.395 -0.845 28.725 -0.515 ;
      RECT 27.715 -1.525 28.045 -1.195 ;
      RECT 27.035 -0.845 27.365 -0.515 ;
      RECT 26.355 -1.525 26.685 -1.195 ;
      RECT 25.675 -0.845 26.005 -0.515 ;
      RECT 24.995 -1.525 25.325 -1.195 ;
      RECT 24.315 -0.845 24.645 -0.515 ;
      RECT 23.635 -1.525 23.965 -1.195 ;
      RECT 22.955 -0.845 23.285 -0.515 ;
      RECT 22.275 -1.525 22.605 -1.195 ;
      RECT 21.595 -0.845 21.925 -0.515 ;
      RECT 20.915 -1.525 21.245 -1.195 ;
      RECT 20.235 -0.845 20.565 -0.515 ;
      RECT 19.555 -1.525 19.885 -1.195 ;
      RECT 18.875 -0.845 19.205 -0.515 ;
      RECT 18.195 -1.525 18.525 -1.195 ;
      RECT 17.515 -0.845 17.845 -0.515 ;
      RECT 16.835 -1.525 17.165 -1.195 ;
      RECT 16.155 -0.845 16.485 -0.515 ;
      RECT 15.475 -1.525 15.805 -1.195 ;
      RECT 14.795 -0.845 15.125 -0.515 ;
      RECT 14.115 -1.525 14.445 -1.195 ;
      RECT 13.435 -0.845 13.765 -0.515 ;
      RECT 12.755 -1.525 13.085 -1.195 ;
      RECT 12.075 -0.845 12.405 -0.515 ;
      RECT 11.395 -1.525 11.725 -1.195 ;
      RECT 10.715 -0.845 11.045 -0.515 ;
      RECT 10.035 -1.525 10.365 -1.195 ;
      RECT 9.355 -0.845 9.685 -0.515 ;
      RECT 8.675 -1.525 9.005 -1.195 ;
      RECT 7.995 -0.845 8.325 -0.515 ;
      RECT 7.315 -1.525 7.645 -1.195 ;
      RECT 6.635 -0.845 6.965 -0.515 ;
      RECT 5.955 -1.525 6.285 -1.195 ;
      RECT 5.275 -0.845 5.605 -0.515 ;
      RECT 4.595 -1.525 4.925 -1.195 ;
      RECT 3.915 -0.845 4.245 -0.515 ;
      RECT 3.235 -1.525 3.565 -1.195 ;
      RECT 2.555 -0.845 2.885 -0.515 ;
      RECT 1.875 -1.525 2.205 -1.195 ;
      RECT 1.195 -0.845 1.525 -0.515 ;
      RECT 0.515 -1.525 0.845 -1.195 ;
      RECT -0.165 -0.845 0.165 -0.515 ;
      RECT -0.845 -1.525 -0.515 -1.195 ;
      RECT -1.525 -0.845 -1.195 -0.515 ;
      RECT -2.205 -1.525 -1.875 -1.195 ;
      RECT -2.88 -0.16 -2.56 7.64 ;
  END
END tristate_inv_delay_line_128

END LIBRARY
