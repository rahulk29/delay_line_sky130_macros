VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO tristate_inv_delay_line_128
  CLASS BLOCK ;
  ORIGIN 2.905 12 ;
  FOREIGN tristate_inv_delay_line_128 -2.905 -12 ;
  SIZE 772.17 BY 35.965 ;
  SYMMETRY X Y R90 ;
  PIN clk_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT -1.47 -12 -1.15 18.92 ;
    END
  END clk_in
  PIN clk_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.52 -12 1.84 18.92 ;
    END
  END clk_out
  PIN ctl[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.03 -12 0.35 18.92 ;
    END
  END ctl[0]
  PIN ctl[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 600.03 -12 600.35 18.92 ;
    END
  END ctl[100]
  PIN ctl[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 606.03 -12 606.35 18.92 ;
    END
  END ctl[101]
  PIN ctl[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 612.03 -12 612.35 18.92 ;
    END
  END ctl[102]
  PIN ctl[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 618.03 -12 618.35 18.92 ;
    END
  END ctl[103]
  PIN ctl[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 624.03 -12 624.35 18.92 ;
    END
  END ctl[104]
  PIN ctl[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 630.03 -12 630.35 18.92 ;
    END
  END ctl[105]
  PIN ctl[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 636.03 -12 636.35 18.92 ;
    END
  END ctl[106]
  PIN ctl[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 642.03 -12 642.35 18.92 ;
    END
  END ctl[107]
  PIN ctl[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 648.03 -12 648.35 18.92 ;
    END
  END ctl[108]
  PIN ctl[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 654.03 -12 654.35 18.92 ;
    END
  END ctl[109]
  PIN ctl[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 60.03 -12 60.35 18.92 ;
    END
  END ctl[10]
  PIN ctl[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 660.03 -12 660.35 18.92 ;
    END
  END ctl[110]
  PIN ctl[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 666.03 -12 666.35 18.92 ;
    END
  END ctl[111]
  PIN ctl[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 672.03 -12 672.35 18.92 ;
    END
  END ctl[112]
  PIN ctl[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 678.03 -12 678.35 18.92 ;
    END
  END ctl[113]
  PIN ctl[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 684.03 -12 684.35 18.92 ;
    END
  END ctl[114]
  PIN ctl[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 690.03 -12 690.35 18.92 ;
    END
  END ctl[115]
  PIN ctl[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 696.03 -12 696.35 18.92 ;
    END
  END ctl[116]
  PIN ctl[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 702.03 -12 702.35 18.92 ;
    END
  END ctl[117]
  PIN ctl[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 708.03 -12 708.35 18.92 ;
    END
  END ctl[118]
  PIN ctl[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 714.03 -12 714.35 18.92 ;
    END
  END ctl[119]
  PIN ctl[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 66.03 -12 66.35 18.92 ;
    END
  END ctl[11]
  PIN ctl[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 720.03 -12 720.35 18.92 ;
    END
  END ctl[120]
  PIN ctl[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 726.03 -12 726.35 18.92 ;
    END
  END ctl[121]
  PIN ctl[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 732.03 -12 732.35 18.92 ;
    END
  END ctl[122]
  PIN ctl[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 738.03 -12 738.35 18.92 ;
    END
  END ctl[123]
  PIN ctl[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 744.03 -12 744.35 18.92 ;
    END
  END ctl[124]
  PIN ctl[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 750.03 -12 750.35 18.92 ;
    END
  END ctl[125]
  PIN ctl[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 756.03 -12 756.35 18.92 ;
    END
  END ctl[126]
  PIN ctl[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 762.03 -12 762.35 18.92 ;
    END
  END ctl[127]
  PIN ctl[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 72.03 -12 72.35 18.92 ;
    END
  END ctl[12]
  PIN ctl[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 78.03 -12 78.35 18.92 ;
    END
  END ctl[13]
  PIN ctl[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 84.03 -12 84.35 18.92 ;
    END
  END ctl[14]
  PIN ctl[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 90.03 -12 90.35 18.92 ;
    END
  END ctl[15]
  PIN ctl[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 96.03 -12 96.35 18.92 ;
    END
  END ctl[16]
  PIN ctl[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 102.03 -12 102.35 18.92 ;
    END
  END ctl[17]
  PIN ctl[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 108.03 -12 108.35 18.92 ;
    END
  END ctl[18]
  PIN ctl[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 114.03 -12 114.35 18.92 ;
    END
  END ctl[19]
  PIN ctl[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 6.03 -12 6.35 18.92 ;
    END
  END ctl[1]
  PIN ctl[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 120.03 -12 120.35 18.92 ;
    END
  END ctl[20]
  PIN ctl[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 126.03 -12 126.35 18.92 ;
    END
  END ctl[21]
  PIN ctl[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 132.03 -12 132.35 18.92 ;
    END
  END ctl[22]
  PIN ctl[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 138.03 -12 138.35 18.92 ;
    END
  END ctl[23]
  PIN ctl[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 144.03 -12 144.35 18.92 ;
    END
  END ctl[24]
  PIN ctl[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 150.03 -12 150.35 18.92 ;
    END
  END ctl[25]
  PIN ctl[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 156.03 -12 156.35 18.92 ;
    END
  END ctl[26]
  PIN ctl[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 162.03 -12 162.35 18.92 ;
    END
  END ctl[27]
  PIN ctl[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 168.03 -12 168.35 18.92 ;
    END
  END ctl[28]
  PIN ctl[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 174.03 -12 174.35 18.92 ;
    END
  END ctl[29]
  PIN ctl[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 12.03 -12 12.35 18.92 ;
    END
  END ctl[2]
  PIN ctl[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 180.03 -12 180.35 18.92 ;
    END
  END ctl[30]
  PIN ctl[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 186.03 -12 186.35 18.92 ;
    END
  END ctl[31]
  PIN ctl[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 192.03 -12 192.35 18.92 ;
    END
  END ctl[32]
  PIN ctl[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 198.03 -12 198.35 18.92 ;
    END
  END ctl[33]
  PIN ctl[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 204.03 -12 204.35 18.92 ;
    END
  END ctl[34]
  PIN ctl[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 210.03 -12 210.35 18.92 ;
    END
  END ctl[35]
  PIN ctl[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 216.03 -12 216.35 18.92 ;
    END
  END ctl[36]
  PIN ctl[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 222.03 -12 222.35 18.92 ;
    END
  END ctl[37]
  PIN ctl[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 228.03 -12 228.35 18.92 ;
    END
  END ctl[38]
  PIN ctl[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 234.03 -12 234.35 18.92 ;
    END
  END ctl[39]
  PIN ctl[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.03 -12 18.35 18.92 ;
    END
  END ctl[3]
  PIN ctl[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 240.03 -12 240.35 18.92 ;
    END
  END ctl[40]
  PIN ctl[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 246.03 -12 246.35 18.92 ;
    END
  END ctl[41]
  PIN ctl[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 252.03 -12 252.35 18.92 ;
    END
  END ctl[42]
  PIN ctl[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 258.03 -12 258.35 18.92 ;
    END
  END ctl[43]
  PIN ctl[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 264.03 -12 264.35 18.92 ;
    END
  END ctl[44]
  PIN ctl[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 270.03 -12 270.35 18.92 ;
    END
  END ctl[45]
  PIN ctl[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 276.03 -12 276.35 18.92 ;
    END
  END ctl[46]
  PIN ctl[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 282.03 -12 282.35 18.92 ;
    END
  END ctl[47]
  PIN ctl[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 288.03 -12 288.35 18.92 ;
    END
  END ctl[48]
  PIN ctl[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 294.03 -12 294.35 18.92 ;
    END
  END ctl[49]
  PIN ctl[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 24.03 -12 24.35 18.92 ;
    END
  END ctl[4]
  PIN ctl[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 300.03 -12 300.35 18.92 ;
    END
  END ctl[50]
  PIN ctl[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 306.03 -12 306.35 18.92 ;
    END
  END ctl[51]
  PIN ctl[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 312.03 -12 312.35 18.92 ;
    END
  END ctl[52]
  PIN ctl[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 318.03 -12 318.35 18.92 ;
    END
  END ctl[53]
  PIN ctl[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 324.03 -12 324.35 18.92 ;
    END
  END ctl[54]
  PIN ctl[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 330.03 -12 330.35 18.92 ;
    END
  END ctl[55]
  PIN ctl[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 336.03 -12 336.35 18.92 ;
    END
  END ctl[56]
  PIN ctl[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 342.03 -12 342.35 18.92 ;
    END
  END ctl[57]
  PIN ctl[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 348.03 -12 348.35 18.92 ;
    END
  END ctl[58]
  PIN ctl[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 354.03 -12 354.35 18.92 ;
    END
  END ctl[59]
  PIN ctl[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 30.03 -12 30.35 18.92 ;
    END
  END ctl[5]
  PIN ctl[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 360.03 -12 360.35 18.92 ;
    END
  END ctl[60]
  PIN ctl[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 366.03 -12 366.35 18.92 ;
    END
  END ctl[61]
  PIN ctl[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 372.03 -12 372.35 18.92 ;
    END
  END ctl[62]
  PIN ctl[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 378.03 -12 378.35 18.92 ;
    END
  END ctl[63]
  PIN ctl[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 384.03 -12 384.35 18.92 ;
    END
  END ctl[64]
  PIN ctl[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 390.03 -12 390.35 18.92 ;
    END
  END ctl[65]
  PIN ctl[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 396.03 -12 396.35 18.92 ;
    END
  END ctl[66]
  PIN ctl[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 402.03 -12 402.35 18.92 ;
    END
  END ctl[67]
  PIN ctl[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 408.03 -12 408.35 18.92 ;
    END
  END ctl[68]
  PIN ctl[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 414.03 -12 414.35 18.92 ;
    END
  END ctl[69]
  PIN ctl[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 36.03 -12 36.35 18.92 ;
    END
  END ctl[6]
  PIN ctl[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 420.03 -12 420.35 18.92 ;
    END
  END ctl[70]
  PIN ctl[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 426.03 -12 426.35 18.92 ;
    END
  END ctl[71]
  PIN ctl[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 432.03 -12 432.35 18.92 ;
    END
  END ctl[72]
  PIN ctl[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 438.03 -12 438.35 18.92 ;
    END
  END ctl[73]
  PIN ctl[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 444.03 -12 444.35 18.92 ;
    END
  END ctl[74]
  PIN ctl[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 450.03 -12 450.35 18.92 ;
    END
  END ctl[75]
  PIN ctl[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 456.03 -12 456.35 18.92 ;
    END
  END ctl[76]
  PIN ctl[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 462.03 -12 462.35 18.92 ;
    END
  END ctl[77]
  PIN ctl[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 468.03 -12 468.35 18.92 ;
    END
  END ctl[78]
  PIN ctl[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 474.03 -12 474.35 18.92 ;
    END
  END ctl[79]
  PIN ctl[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 42.03 -12 42.35 18.92 ;
    END
  END ctl[7]
  PIN ctl[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 480.03 -12 480.35 18.92 ;
    END
  END ctl[80]
  PIN ctl[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 486.03 -12 486.35 18.92 ;
    END
  END ctl[81]
  PIN ctl[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 492.03 -12 492.35 18.92 ;
    END
  END ctl[82]
  PIN ctl[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 498.03 -12 498.35 18.92 ;
    END
  END ctl[83]
  PIN ctl[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 504.03 -12 504.35 18.92 ;
    END
  END ctl[84]
  PIN ctl[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 510.03 -12 510.35 18.92 ;
    END
  END ctl[85]
  PIN ctl[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 516.03 -12 516.35 18.92 ;
    END
  END ctl[86]
  PIN ctl[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 522.03 -12 522.35 18.92 ;
    END
  END ctl[87]
  PIN ctl[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 528.03 -12 528.35 18.92 ;
    END
  END ctl[88]
  PIN ctl[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 534.03 -12 534.35 18.92 ;
    END
  END ctl[89]
  PIN ctl[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 48.03 -12 48.35 18.92 ;
    END
  END ctl[8]
  PIN ctl[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 540.03 -12 540.35 18.92 ;
    END
  END ctl[90]
  PIN ctl[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 546.03 -12 546.35 18.92 ;
    END
  END ctl[91]
  PIN ctl[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 552.03 -12 552.35 18.92 ;
    END
  END ctl[92]
  PIN ctl[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 558.03 -12 558.35 18.92 ;
    END
  END ctl[93]
  PIN ctl[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 564.03 -12 564.35 18.92 ;
    END
  END ctl[94]
  PIN ctl[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 570.03 -12 570.35 18.92 ;
    END
  END ctl[95]
  PIN ctl[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 576.03 -12 576.35 18.92 ;
    END
  END ctl[96]
  PIN ctl[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 582.03 -12 582.35 18.92 ;
    END
  END ctl[97]
  PIN ctl[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 588.03 -12 588.35 18.92 ;
    END
  END ctl[98]
  PIN ctl[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 594.03 -12 594.35 18.92 ;
    END
  END ctl[99]
  PIN ctl[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 54.03 -12 54.35 18.92 ;
    END
  END ctl[9]
  PIN ctl_b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 4.05 -12 4.37 18.92 ;
    END
  END ctl_b[0]
  PIN ctl_b[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 604.05 -12 604.37 18.92 ;
    END
  END ctl_b[100]
  PIN ctl_b[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 610.05 -12 610.37 18.92 ;
    END
  END ctl_b[101]
  PIN ctl_b[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 616.05 -12 616.37 18.92 ;
    END
  END ctl_b[102]
  PIN ctl_b[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 622.05 -12 622.37 18.92 ;
    END
  END ctl_b[103]
  PIN ctl_b[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 628.05 -12 628.37 18.92 ;
    END
  END ctl_b[104]
  PIN ctl_b[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 634.05 -12 634.37 18.92 ;
    END
  END ctl_b[105]
  PIN ctl_b[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 640.05 -12 640.37 18.92 ;
    END
  END ctl_b[106]
  PIN ctl_b[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 646.05 -12 646.37 18.92 ;
    END
  END ctl_b[107]
  PIN ctl_b[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 652.05 -12 652.37 18.92 ;
    END
  END ctl_b[108]
  PIN ctl_b[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 658.05 -12 658.37 18.92 ;
    END
  END ctl_b[109]
  PIN ctl_b[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 64.05 -12 64.37 18.92 ;
    END
  END ctl_b[10]
  PIN ctl_b[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 664.05 -12 664.37 18.92 ;
    END
  END ctl_b[110]
  PIN ctl_b[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 670.05 -12 670.37 18.92 ;
    END
  END ctl_b[111]
  PIN ctl_b[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 676.05 -12 676.37 18.92 ;
    END
  END ctl_b[112]
  PIN ctl_b[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 682.05 -12 682.37 18.92 ;
    END
  END ctl_b[113]
  PIN ctl_b[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 688.05 -12 688.37 18.92 ;
    END
  END ctl_b[114]
  PIN ctl_b[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 694.05 -12 694.37 18.92 ;
    END
  END ctl_b[115]
  PIN ctl_b[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 700.05 -12 700.37 18.92 ;
    END
  END ctl_b[116]
  PIN ctl_b[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 706.05 -12 706.37 18.92 ;
    END
  END ctl_b[117]
  PIN ctl_b[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 712.05 -12 712.37 18.92 ;
    END
  END ctl_b[118]
  PIN ctl_b[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 718.05 -12 718.37 18.92 ;
    END
  END ctl_b[119]
  PIN ctl_b[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 70.05 -12 70.37 18.92 ;
    END
  END ctl_b[11]
  PIN ctl_b[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 724.05 -12 724.37 18.92 ;
    END
  END ctl_b[120]
  PIN ctl_b[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 730.05 -12 730.37 18.92 ;
    END
  END ctl_b[121]
  PIN ctl_b[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 736.05 -12 736.37 18.92 ;
    END
  END ctl_b[122]
  PIN ctl_b[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 742.05 -12 742.37 18.92 ;
    END
  END ctl_b[123]
  PIN ctl_b[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 748.05 -12 748.37 18.92 ;
    END
  END ctl_b[124]
  PIN ctl_b[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 754.05 -12 754.37 18.92 ;
    END
  END ctl_b[125]
  PIN ctl_b[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 760.05 -12 760.37 18.92 ;
    END
  END ctl_b[126]
  PIN ctl_b[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 766.05 -12 766.37 18.92 ;
    END
  END ctl_b[127]
  PIN ctl_b[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 76.05 -12 76.37 18.92 ;
    END
  END ctl_b[12]
  PIN ctl_b[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 82.05 -12 82.37 18.92 ;
    END
  END ctl_b[13]
  PIN ctl_b[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 88.05 -12 88.37 18.92 ;
    END
  END ctl_b[14]
  PIN ctl_b[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 94.05 -12 94.37 18.92 ;
    END
  END ctl_b[15]
  PIN ctl_b[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 100.05 -12 100.37 18.92 ;
    END
  END ctl_b[16]
  PIN ctl_b[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 106.05 -12 106.37 18.92 ;
    END
  END ctl_b[17]
  PIN ctl_b[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 112.05 -12 112.37 18.92 ;
    END
  END ctl_b[18]
  PIN ctl_b[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 118.05 -12 118.37 18.92 ;
    END
  END ctl_b[19]
  PIN ctl_b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 10.05 -12 10.37 18.92 ;
    END
  END ctl_b[1]
  PIN ctl_b[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 124.05 -12 124.37 18.92 ;
    END
  END ctl_b[20]
  PIN ctl_b[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 130.05 -12 130.37 18.92 ;
    END
  END ctl_b[21]
  PIN ctl_b[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 136.05 -12 136.37 18.92 ;
    END
  END ctl_b[22]
  PIN ctl_b[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 142.05 -12 142.37 18.92 ;
    END
  END ctl_b[23]
  PIN ctl_b[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 148.05 -12 148.37 18.92 ;
    END
  END ctl_b[24]
  PIN ctl_b[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 154.05 -12 154.37 18.92 ;
    END
  END ctl_b[25]
  PIN ctl_b[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 160.05 -12 160.37 18.92 ;
    END
  END ctl_b[26]
  PIN ctl_b[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 166.05 -12 166.37 18.92 ;
    END
  END ctl_b[27]
  PIN ctl_b[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 172.05 -12 172.37 18.92 ;
    END
  END ctl_b[28]
  PIN ctl_b[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 178.05 -12 178.37 18.92 ;
    END
  END ctl_b[29]
  PIN ctl_b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.05 -12 16.37 18.92 ;
    END
  END ctl_b[2]
  PIN ctl_b[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 184.05 -12 184.37 18.92 ;
    END
  END ctl_b[30]
  PIN ctl_b[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 190.05 -12 190.37 18.92 ;
    END
  END ctl_b[31]
  PIN ctl_b[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 196.05 -12 196.37 18.92 ;
    END
  END ctl_b[32]
  PIN ctl_b[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 202.05 -12 202.37 18.92 ;
    END
  END ctl_b[33]
  PIN ctl_b[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 208.05 -12 208.37 18.92 ;
    END
  END ctl_b[34]
  PIN ctl_b[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 214.05 -12 214.37 18.92 ;
    END
  END ctl_b[35]
  PIN ctl_b[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 220.05 -12 220.37 18.92 ;
    END
  END ctl_b[36]
  PIN ctl_b[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 226.05 -12 226.37 18.92 ;
    END
  END ctl_b[37]
  PIN ctl_b[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 232.05 -12 232.37 18.92 ;
    END
  END ctl_b[38]
  PIN ctl_b[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 238.05 -12 238.37 18.92 ;
    END
  END ctl_b[39]
  PIN ctl_b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 22.05 -12 22.37 18.92 ;
    END
  END ctl_b[3]
  PIN ctl_b[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 244.05 -12 244.37 18.92 ;
    END
  END ctl_b[40]
  PIN ctl_b[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 250.05 -12 250.37 18.92 ;
    END
  END ctl_b[41]
  PIN ctl_b[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 256.05 -12 256.37 18.92 ;
    END
  END ctl_b[42]
  PIN ctl_b[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 262.05 -12 262.37 18.92 ;
    END
  END ctl_b[43]
  PIN ctl_b[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 268.05 -12 268.37 18.92 ;
    END
  END ctl_b[44]
  PIN ctl_b[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 274.05 -12 274.37 18.92 ;
    END
  END ctl_b[45]
  PIN ctl_b[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 280.05 -12 280.37 18.92 ;
    END
  END ctl_b[46]
  PIN ctl_b[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 286.05 -12 286.37 18.92 ;
    END
  END ctl_b[47]
  PIN ctl_b[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 292.05 -12 292.37 18.92 ;
    END
  END ctl_b[48]
  PIN ctl_b[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 298.05 -12 298.37 18.92 ;
    END
  END ctl_b[49]
  PIN ctl_b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 28.05 -12 28.37 18.92 ;
    END
  END ctl_b[4]
  PIN ctl_b[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 304.05 -12 304.37 18.92 ;
    END
  END ctl_b[50]
  PIN ctl_b[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 310.05 -12 310.37 18.92 ;
    END
  END ctl_b[51]
  PIN ctl_b[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 316.05 -12 316.37 18.92 ;
    END
  END ctl_b[52]
  PIN ctl_b[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 322.05 -12 322.37 18.92 ;
    END
  END ctl_b[53]
  PIN ctl_b[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 328.05 -12 328.37 18.92 ;
    END
  END ctl_b[54]
  PIN ctl_b[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 334.05 -12 334.37 18.92 ;
    END
  END ctl_b[55]
  PIN ctl_b[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 340.05 -12 340.37 18.92 ;
    END
  END ctl_b[56]
  PIN ctl_b[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 346.05 -12 346.37 18.92 ;
    END
  END ctl_b[57]
  PIN ctl_b[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 352.05 -12 352.37 18.92 ;
    END
  END ctl_b[58]
  PIN ctl_b[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 358.05 -12 358.37 18.92 ;
    END
  END ctl_b[59]
  PIN ctl_b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 34.05 -12 34.37 18.92 ;
    END
  END ctl_b[5]
  PIN ctl_b[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 364.05 -12 364.37 18.92 ;
    END
  END ctl_b[60]
  PIN ctl_b[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 370.05 -12 370.37 18.92 ;
    END
  END ctl_b[61]
  PIN ctl_b[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 376.05 -12 376.37 18.92 ;
    END
  END ctl_b[62]
  PIN ctl_b[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 382.05 -12 382.37 18.92 ;
    END
  END ctl_b[63]
  PIN ctl_b[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 388.05 -12 388.37 18.92 ;
    END
  END ctl_b[64]
  PIN ctl_b[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 394.05 -12 394.37 18.92 ;
    END
  END ctl_b[65]
  PIN ctl_b[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 400.05 -12 400.37 18.92 ;
    END
  END ctl_b[66]
  PIN ctl_b[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 406.05 -12 406.37 18.92 ;
    END
  END ctl_b[67]
  PIN ctl_b[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 412.05 -12 412.37 18.92 ;
    END
  END ctl_b[68]
  PIN ctl_b[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 418.05 -12 418.37 18.92 ;
    END
  END ctl_b[69]
  PIN ctl_b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 40.05 -12 40.37 18.92 ;
    END
  END ctl_b[6]
  PIN ctl_b[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 424.05 -12 424.37 18.92 ;
    END
  END ctl_b[70]
  PIN ctl_b[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 430.05 -12 430.37 18.92 ;
    END
  END ctl_b[71]
  PIN ctl_b[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 436.05 -12 436.37 18.92 ;
    END
  END ctl_b[72]
  PIN ctl_b[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 442.05 -12 442.37 18.92 ;
    END
  END ctl_b[73]
  PIN ctl_b[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 448.05 -12 448.37 18.92 ;
    END
  END ctl_b[74]
  PIN ctl_b[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 454.05 -12 454.37 18.92 ;
    END
  END ctl_b[75]
  PIN ctl_b[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 460.05 -12 460.37 18.92 ;
    END
  END ctl_b[76]
  PIN ctl_b[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 466.05 -12 466.37 18.92 ;
    END
  END ctl_b[77]
  PIN ctl_b[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 472.05 -12 472.37 18.92 ;
    END
  END ctl_b[78]
  PIN ctl_b[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 478.05 -12 478.37 18.92 ;
    END
  END ctl_b[79]
  PIN ctl_b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 46.05 -12 46.37 18.92 ;
    END
  END ctl_b[7]
  PIN ctl_b[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 484.05 -12 484.37 18.92 ;
    END
  END ctl_b[80]
  PIN ctl_b[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 490.05 -12 490.37 18.92 ;
    END
  END ctl_b[81]
  PIN ctl_b[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 496.05 -12 496.37 18.92 ;
    END
  END ctl_b[82]
  PIN ctl_b[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 502.05 -12 502.37 18.92 ;
    END
  END ctl_b[83]
  PIN ctl_b[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 508.05 -12 508.37 18.92 ;
    END
  END ctl_b[84]
  PIN ctl_b[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 514.05 -12 514.37 18.92 ;
    END
  END ctl_b[85]
  PIN ctl_b[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 520.05 -12 520.37 18.92 ;
    END
  END ctl_b[86]
  PIN ctl_b[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 526.05 -12 526.37 18.92 ;
    END
  END ctl_b[87]
  PIN ctl_b[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 532.05 -12 532.37 18.92 ;
    END
  END ctl_b[88]
  PIN ctl_b[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 538.05 -12 538.37 18.92 ;
    END
  END ctl_b[89]
  PIN ctl_b[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 52.05 -12 52.37 18.92 ;
    END
  END ctl_b[8]
  PIN ctl_b[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 544.05 -12 544.37 18.92 ;
    END
  END ctl_b[90]
  PIN ctl_b[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 550.05 -12 550.37 18.92 ;
    END
  END ctl_b[91]
  PIN ctl_b[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 556.05 -12 556.37 18.92 ;
    END
  END ctl_b[92]
  PIN ctl_b[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 562.05 -12 562.37 18.92 ;
    END
  END ctl_b[93]
  PIN ctl_b[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 568.05 -12 568.37 18.92 ;
    END
  END ctl_b[94]
  PIN ctl_b[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 574.05 -12 574.37 18.92 ;
    END
  END ctl_b[95]
  PIN ctl_b[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 580.05 -12 580.37 18.92 ;
    END
  END ctl_b[96]
  PIN ctl_b[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 586.05 -12 586.37 18.92 ;
    END
  END ctl_b[97]
  PIN ctl_b[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 592.05 -12 592.37 18.92 ;
    END
  END ctl_b[98]
  PIN ctl_b[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 598.05 -12 598.37 18.92 ;
    END
  END ctl_b[99]
  PIN ctl_b[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 58.05 -12 58.37 18.92 ;
    END
  END ctl_b[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 641.075 15.475 641.405 15.805 ;
        RECT 641.075 11.395 641.405 11.725 ;
        RECT 641.075 10.035 641.405 10.365 ;
        RECT 641.075 8.675 641.405 9.005 ;
        RECT 641.075 7.315 641.405 7.645 ;
        RECT 641.075 5.955 641.405 6.285 ;
        RECT 641.075 4.595 641.405 4.925 ;
        RECT 641.075 3.235 641.405 3.565 ;
        RECT 641.075 1.875 641.405 2.205 ;
        RECT 641.075 0.515 641.405 0.845 ;
        RECT 641.08 -8.32 641.4 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 642.435 15.475 642.765 15.805 ;
        RECT 642.435 11.395 642.765 11.725 ;
        RECT 642.435 10.035 642.765 10.365 ;
        RECT 642.435 8.675 642.765 9.005 ;
        RECT 642.435 7.315 642.765 7.645 ;
        RECT 642.435 5.955 642.765 6.285 ;
        RECT 642.435 4.595 642.765 4.925 ;
        RECT 642.435 3.235 642.765 3.565 ;
        RECT 642.435 1.875 642.765 2.205 ;
        RECT 642.435 0.515 642.765 0.845 ;
        RECT 642.44 -8.32 642.76 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 643.795 15.475 644.125 15.805 ;
        RECT 643.795 10.035 644.125 10.365 ;
        RECT 643.795 8.675 644.125 9.005 ;
        RECT 643.795 7.315 644.125 7.645 ;
        RECT 643.795 5.955 644.125 6.285 ;
        RECT 643.795 4.595 644.125 4.925 ;
        RECT 643.795 3.235 644.125 3.565 ;
        RECT 643.795 1.875 644.125 2.205 ;
        RECT 643.795 0.515 644.125 0.845 ;
        RECT 643.8 -8.32 644.12 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 645.155 15.475 645.485 15.805 ;
        RECT 645.155 10.035 645.485 10.365 ;
        RECT 645.155 8.675 645.485 9.005 ;
        RECT 645.155 7.315 645.485 7.645 ;
        RECT 645.155 5.955 645.485 6.285 ;
        RECT 645.155 4.595 645.485 4.925 ;
        RECT 645.155 3.235 645.485 3.565 ;
        RECT 645.155 1.875 645.485 2.205 ;
        RECT 645.155 0.515 645.485 0.845 ;
        RECT 645.16 -8.32 645.48 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 646.515 15.475 646.845 15.805 ;
        RECT 646.515 10.035 646.845 10.365 ;
        RECT 646.515 8.675 646.845 9.005 ;
        RECT 646.515 7.315 646.845 7.645 ;
        RECT 646.515 5.955 646.845 6.285 ;
        RECT 646.515 4.595 646.845 4.925 ;
        RECT 646.515 3.235 646.845 3.565 ;
        RECT 646.515 1.875 646.845 2.205 ;
        RECT 646.515 0.515 646.845 0.845 ;
        RECT 646.52 -8.32 646.84 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 647.875 15.475 648.205 15.805 ;
        RECT 647.875 10.035 648.205 10.365 ;
        RECT 647.875 8.675 648.205 9.005 ;
        RECT 647.875 7.315 648.205 7.645 ;
        RECT 647.875 5.955 648.205 6.285 ;
        RECT 647.875 4.595 648.205 4.925 ;
        RECT 647.875 3.235 648.205 3.565 ;
        RECT 647.875 1.875 648.205 2.205 ;
        RECT 647.875 0.515 648.205 0.845 ;
        RECT 647.88 -8.32 648.2 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 649.235 15.475 649.565 15.805 ;
        RECT 649.235 10.035 649.565 10.365 ;
        RECT 649.235 8.675 649.565 9.005 ;
        RECT 649.235 7.315 649.565 7.645 ;
        RECT 649.235 5.955 649.565 6.285 ;
        RECT 649.235 4.595 649.565 4.925 ;
        RECT 649.235 3.235 649.565 3.565 ;
        RECT 649.235 1.875 649.565 2.205 ;
        RECT 649.235 0.515 649.565 0.845 ;
        RECT 649.24 -8.32 649.56 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 650.595 15.475 650.925 15.805 ;
        RECT 650.595 10.035 650.925 10.365 ;
        RECT 650.595 8.675 650.925 9.005 ;
        RECT 650.595 7.315 650.925 7.645 ;
        RECT 650.595 5.955 650.925 6.285 ;
        RECT 650.595 4.595 650.925 4.925 ;
        RECT 650.595 3.235 650.925 3.565 ;
        RECT 650.595 1.875 650.925 2.205 ;
        RECT 650.595 0.515 650.925 0.845 ;
        RECT 650.6 -8.32 650.92 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 651.955 15.475 652.285 15.805 ;
        RECT 651.955 11.395 652.285 11.725 ;
        RECT 651.955 10.035 652.285 10.365 ;
        RECT 651.955 8.675 652.285 9.005 ;
        RECT 651.955 7.315 652.285 7.645 ;
        RECT 651.955 5.955 652.285 6.285 ;
        RECT 651.955 4.595 652.285 4.925 ;
        RECT 651.955 3.235 652.285 3.565 ;
        RECT 651.955 1.875 652.285 2.205 ;
        RECT 651.955 0.515 652.285 0.845 ;
        RECT 651.96 -8.32 652.28 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 653.315 15.475 653.645 15.805 ;
        RECT 653.315 11.395 653.645 11.725 ;
        RECT 653.315 10.035 653.645 10.365 ;
        RECT 653.315 8.675 653.645 9.005 ;
        RECT 653.315 7.315 653.645 7.645 ;
        RECT 653.315 5.955 653.645 6.285 ;
        RECT 653.315 4.595 653.645 4.925 ;
        RECT 653.315 3.235 653.645 3.565 ;
        RECT 653.315 1.875 653.645 2.205 ;
        RECT 653.315 0.515 653.645 0.845 ;
        RECT 653.32 -8.32 653.64 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 654.675 15.475 655.005 15.805 ;
        RECT 654.675 11.395 655.005 11.725 ;
        RECT 654.675 10.035 655.005 10.365 ;
        RECT 654.675 8.675 655.005 9.005 ;
        RECT 654.675 7.315 655.005 7.645 ;
        RECT 654.675 5.955 655.005 6.285 ;
        RECT 654.675 4.595 655.005 4.925 ;
        RECT 654.675 3.235 655.005 3.565 ;
        RECT 654.675 1.875 655.005 2.205 ;
        RECT 654.675 0.515 655.005 0.845 ;
        RECT 654.68 -8.32 655 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 656.035 15.475 656.365 15.805 ;
        RECT 656.035 10.035 656.365 10.365 ;
        RECT 656.035 8.675 656.365 9.005 ;
        RECT 656.035 7.315 656.365 7.645 ;
        RECT 656.035 5.955 656.365 6.285 ;
        RECT 656.035 4.595 656.365 4.925 ;
        RECT 656.035 3.235 656.365 3.565 ;
        RECT 656.035 1.875 656.365 2.205 ;
        RECT 656.035 0.515 656.365 0.845 ;
        RECT 656.04 -8.32 656.36 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 657.395 15.475 657.725 15.805 ;
        RECT 657.395 10.035 657.725 10.365 ;
        RECT 657.395 8.675 657.725 9.005 ;
        RECT 657.395 7.315 657.725 7.645 ;
        RECT 657.395 5.955 657.725 6.285 ;
        RECT 657.395 4.595 657.725 4.925 ;
        RECT 657.395 3.235 657.725 3.565 ;
        RECT 657.395 1.875 657.725 2.205 ;
        RECT 657.395 0.515 657.725 0.845 ;
        RECT 657.4 -8.32 657.72 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 658.755 15.475 659.085 15.805 ;
        RECT 658.755 10.035 659.085 10.365 ;
        RECT 658.755 8.675 659.085 9.005 ;
        RECT 658.755 7.315 659.085 7.645 ;
        RECT 658.755 5.955 659.085 6.285 ;
        RECT 658.755 4.595 659.085 4.925 ;
        RECT 658.755 3.235 659.085 3.565 ;
        RECT 658.755 1.875 659.085 2.205 ;
        RECT 658.755 0.515 659.085 0.845 ;
        RECT 658.76 -8.32 659.08 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 660.115 15.475 660.445 15.805 ;
        RECT 660.115 10.035 660.445 10.365 ;
        RECT 660.115 8.675 660.445 9.005 ;
        RECT 660.115 7.315 660.445 7.645 ;
        RECT 660.115 5.955 660.445 6.285 ;
        RECT 660.115 4.595 660.445 4.925 ;
        RECT 660.115 3.235 660.445 3.565 ;
        RECT 660.115 1.875 660.445 2.205 ;
        RECT 660.115 0.515 660.445 0.845 ;
        RECT 660.12 -8.32 660.44 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 661.475 15.475 661.805 15.805 ;
        RECT 661.475 10.035 661.805 10.365 ;
        RECT 661.475 8.675 661.805 9.005 ;
        RECT 661.475 7.315 661.805 7.645 ;
        RECT 661.475 5.955 661.805 6.285 ;
        RECT 661.475 4.595 661.805 4.925 ;
        RECT 661.475 3.235 661.805 3.565 ;
        RECT 661.475 1.875 661.805 2.205 ;
        RECT 661.475 0.515 661.805 0.845 ;
        RECT 661.48 -8.32 661.8 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 662.835 15.475 663.165 15.805 ;
        RECT 662.835 11.395 663.165 11.725 ;
        RECT 662.835 10.035 663.165 10.365 ;
        RECT 662.835 8.675 663.165 9.005 ;
        RECT 662.835 7.315 663.165 7.645 ;
        RECT 662.835 5.955 663.165 6.285 ;
        RECT 662.835 4.595 663.165 4.925 ;
        RECT 662.835 3.235 663.165 3.565 ;
        RECT 662.835 1.875 663.165 2.205 ;
        RECT 662.835 0.515 663.165 0.845 ;
        RECT 662.84 -8.32 663.16 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 664.195 15.475 664.525 15.805 ;
        RECT 664.195 11.395 664.525 11.725 ;
        RECT 664.195 10.035 664.525 10.365 ;
        RECT 664.195 8.675 664.525 9.005 ;
        RECT 664.195 7.315 664.525 7.645 ;
        RECT 664.195 5.955 664.525 6.285 ;
        RECT 664.195 4.595 664.525 4.925 ;
        RECT 664.195 3.235 664.525 3.565 ;
        RECT 664.195 1.875 664.525 2.205 ;
        RECT 664.195 0.515 664.525 0.845 ;
        RECT 664.2 -8.32 664.52 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 665.555 15.475 665.885 15.805 ;
        RECT 665.555 11.395 665.885 11.725 ;
        RECT 665.555 10.035 665.885 10.365 ;
        RECT 665.555 8.675 665.885 9.005 ;
        RECT 665.555 7.315 665.885 7.645 ;
        RECT 665.555 5.955 665.885 6.285 ;
        RECT 665.555 4.595 665.885 4.925 ;
        RECT 665.555 3.235 665.885 3.565 ;
        RECT 665.555 1.875 665.885 2.205 ;
        RECT 665.555 0.515 665.885 0.845 ;
        RECT 665.56 -8.32 665.88 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 666.915 15.475 667.245 15.805 ;
        RECT 666.915 10.035 667.245 10.365 ;
        RECT 666.915 8.675 667.245 9.005 ;
        RECT 666.915 7.315 667.245 7.645 ;
        RECT 666.915 5.955 667.245 6.285 ;
        RECT 666.915 4.595 667.245 4.925 ;
        RECT 666.915 3.235 667.245 3.565 ;
        RECT 666.915 1.875 667.245 2.205 ;
        RECT 666.915 0.515 667.245 0.845 ;
        RECT 666.92 -8.32 667.24 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 668.275 15.475 668.605 15.805 ;
        RECT 668.275 10.035 668.605 10.365 ;
        RECT 668.275 8.675 668.605 9.005 ;
        RECT 668.275 7.315 668.605 7.645 ;
        RECT 668.275 5.955 668.605 6.285 ;
        RECT 668.275 4.595 668.605 4.925 ;
        RECT 668.275 3.235 668.605 3.565 ;
        RECT 668.275 1.875 668.605 2.205 ;
        RECT 668.275 0.515 668.605 0.845 ;
        RECT 668.28 -8.32 668.6 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 669.635 15.475 669.965 15.805 ;
        RECT 669.635 10.035 669.965 10.365 ;
        RECT 669.635 8.675 669.965 9.005 ;
        RECT 669.635 7.315 669.965 7.645 ;
        RECT 669.635 5.955 669.965 6.285 ;
        RECT 669.635 4.595 669.965 4.925 ;
        RECT 669.635 3.235 669.965 3.565 ;
        RECT 669.635 1.875 669.965 2.205 ;
        RECT 669.635 0.515 669.965 0.845 ;
        RECT 669.64 -8.32 669.96 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 670.995 15.475 671.325 15.805 ;
        RECT 670.995 10.035 671.325 10.365 ;
        RECT 670.995 8.675 671.325 9.005 ;
        RECT 670.995 7.315 671.325 7.645 ;
        RECT 670.995 5.955 671.325 6.285 ;
        RECT 670.995 4.595 671.325 4.925 ;
        RECT 670.995 3.235 671.325 3.565 ;
        RECT 670.995 1.875 671.325 2.205 ;
        RECT 670.995 0.515 671.325 0.845 ;
        RECT 671 -8.32 671.32 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 672.355 15.475 672.685 15.805 ;
        RECT 672.355 10.035 672.685 10.365 ;
        RECT 672.355 8.675 672.685 9.005 ;
        RECT 672.355 7.315 672.685 7.645 ;
        RECT 672.355 5.955 672.685 6.285 ;
        RECT 672.355 4.595 672.685 4.925 ;
        RECT 672.355 3.235 672.685 3.565 ;
        RECT 672.355 1.875 672.685 2.205 ;
        RECT 672.355 0.515 672.685 0.845 ;
        RECT 672.36 -8.32 672.68 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 673.715 15.475 674.045 15.805 ;
        RECT 673.715 10.035 674.045 10.365 ;
        RECT 673.715 8.675 674.045 9.005 ;
        RECT 673.715 7.315 674.045 7.645 ;
        RECT 673.715 5.955 674.045 6.285 ;
        RECT 673.715 4.595 674.045 4.925 ;
        RECT 673.715 3.235 674.045 3.565 ;
        RECT 673.715 1.875 674.045 2.205 ;
        RECT 673.715 0.515 674.045 0.845 ;
        RECT 673.72 -8.32 674.04 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 675.075 15.475 675.405 15.805 ;
        RECT 675.075 11.395 675.405 11.725 ;
        RECT 675.075 10.035 675.405 10.365 ;
        RECT 675.075 8.675 675.405 9.005 ;
        RECT 675.075 7.315 675.405 7.645 ;
        RECT 675.075 5.955 675.405 6.285 ;
        RECT 675.075 4.595 675.405 4.925 ;
        RECT 675.075 3.235 675.405 3.565 ;
        RECT 675.075 1.875 675.405 2.205 ;
        RECT 675.075 0.515 675.405 0.845 ;
        RECT 675.08 -8.32 675.4 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 676.435 15.475 676.765 15.805 ;
        RECT 676.435 11.395 676.765 11.725 ;
        RECT 676.435 10.035 676.765 10.365 ;
        RECT 676.435 8.675 676.765 9.005 ;
        RECT 676.435 7.315 676.765 7.645 ;
        RECT 676.435 5.955 676.765 6.285 ;
        RECT 676.435 4.595 676.765 4.925 ;
        RECT 676.435 3.235 676.765 3.565 ;
        RECT 676.435 1.875 676.765 2.205 ;
        RECT 676.435 0.515 676.765 0.845 ;
        RECT 676.44 -8.32 676.76 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 677.795 15.475 678.125 15.805 ;
        RECT 677.795 11.395 678.125 11.725 ;
        RECT 677.795 10.035 678.125 10.365 ;
        RECT 677.795 8.675 678.125 9.005 ;
        RECT 677.795 7.315 678.125 7.645 ;
        RECT 677.795 5.955 678.125 6.285 ;
        RECT 677.795 4.595 678.125 4.925 ;
        RECT 677.795 3.235 678.125 3.565 ;
        RECT 677.795 1.875 678.125 2.205 ;
        RECT 677.795 0.515 678.125 0.845 ;
        RECT 677.8 -8.32 678.12 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 679.155 15.475 679.485 15.805 ;
        RECT 679.155 10.035 679.485 10.365 ;
        RECT 679.155 8.675 679.485 9.005 ;
        RECT 679.155 7.315 679.485 7.645 ;
        RECT 679.155 5.955 679.485 6.285 ;
        RECT 679.155 4.595 679.485 4.925 ;
        RECT 679.155 3.235 679.485 3.565 ;
        RECT 679.155 1.875 679.485 2.205 ;
        RECT 679.155 0.515 679.485 0.845 ;
        RECT 679.16 -8.32 679.48 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 680.515 15.475 680.845 15.805 ;
        RECT 680.515 10.035 680.845 10.365 ;
        RECT 680.515 8.675 680.845 9.005 ;
        RECT 680.515 7.315 680.845 7.645 ;
        RECT 680.515 5.955 680.845 6.285 ;
        RECT 680.515 4.595 680.845 4.925 ;
        RECT 680.515 3.235 680.845 3.565 ;
        RECT 680.515 1.875 680.845 2.205 ;
        RECT 680.515 0.515 680.845 0.845 ;
        RECT 680.52 -8.32 680.84 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 681.875 15.475 682.205 15.805 ;
        RECT 681.875 10.035 682.205 10.365 ;
        RECT 681.875 8.675 682.205 9.005 ;
        RECT 681.875 7.315 682.205 7.645 ;
        RECT 681.875 5.955 682.205 6.285 ;
        RECT 681.875 4.595 682.205 4.925 ;
        RECT 681.875 3.235 682.205 3.565 ;
        RECT 681.875 1.875 682.205 2.205 ;
        RECT 681.875 0.515 682.205 0.845 ;
        RECT 681.88 -8.32 682.2 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 683.235 15.475 683.565 15.805 ;
        RECT 683.235 10.035 683.565 10.365 ;
        RECT 683.235 8.675 683.565 9.005 ;
        RECT 683.235 7.315 683.565 7.645 ;
        RECT 683.235 5.955 683.565 6.285 ;
        RECT 683.235 4.595 683.565 4.925 ;
        RECT 683.235 3.235 683.565 3.565 ;
        RECT 683.235 1.875 683.565 2.205 ;
        RECT 683.235 0.515 683.565 0.845 ;
        RECT 683.24 -8.32 683.56 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 684.595 15.475 684.925 15.805 ;
        RECT 684.595 10.035 684.925 10.365 ;
        RECT 684.595 8.675 684.925 9.005 ;
        RECT 684.595 7.315 684.925 7.645 ;
        RECT 684.595 5.955 684.925 6.285 ;
        RECT 684.595 4.595 684.925 4.925 ;
        RECT 684.595 3.235 684.925 3.565 ;
        RECT 684.595 1.875 684.925 2.205 ;
        RECT 684.595 0.515 684.925 0.845 ;
        RECT 684.6 -8.32 684.92 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 685.955 15.475 686.285 15.805 ;
        RECT 685.955 10.035 686.285 10.365 ;
        RECT 685.955 8.675 686.285 9.005 ;
        RECT 685.955 7.315 686.285 7.645 ;
        RECT 685.955 5.955 686.285 6.285 ;
        RECT 685.955 4.595 686.285 4.925 ;
        RECT 685.955 3.235 686.285 3.565 ;
        RECT 685.955 1.875 686.285 2.205 ;
        RECT 685.955 0.515 686.285 0.845 ;
        RECT 685.96 -8.32 686.28 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 687.315 15.475 687.645 15.805 ;
        RECT 687.315 11.395 687.645 11.725 ;
        RECT 687.315 10.035 687.645 10.365 ;
        RECT 687.315 8.675 687.645 9.005 ;
        RECT 687.315 7.315 687.645 7.645 ;
        RECT 687.315 5.955 687.645 6.285 ;
        RECT 687.315 4.595 687.645 4.925 ;
        RECT 687.315 3.235 687.645 3.565 ;
        RECT 687.315 1.875 687.645 2.205 ;
        RECT 687.315 0.515 687.645 0.845 ;
        RECT 687.32 -8.32 687.64 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 688.675 15.475 689.005 15.805 ;
        RECT 688.675 11.395 689.005 11.725 ;
        RECT 688.675 10.035 689.005 10.365 ;
        RECT 688.675 8.675 689.005 9.005 ;
        RECT 688.675 7.315 689.005 7.645 ;
        RECT 688.675 5.955 689.005 6.285 ;
        RECT 688.675 4.595 689.005 4.925 ;
        RECT 688.675 3.235 689.005 3.565 ;
        RECT 688.675 1.875 689.005 2.205 ;
        RECT 688.675 0.515 689.005 0.845 ;
        RECT 688.68 -8.32 689 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 690.035 15.475 690.365 15.805 ;
        RECT 690.035 11.395 690.365 11.725 ;
        RECT 690.035 10.035 690.365 10.365 ;
        RECT 690.035 8.675 690.365 9.005 ;
        RECT 690.035 7.315 690.365 7.645 ;
        RECT 690.035 5.955 690.365 6.285 ;
        RECT 690.035 4.595 690.365 4.925 ;
        RECT 690.035 3.235 690.365 3.565 ;
        RECT 690.035 1.875 690.365 2.205 ;
        RECT 690.035 0.515 690.365 0.845 ;
        RECT 690.04 -8.32 690.36 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 691.395 15.475 691.725 15.805 ;
        RECT 691.395 10.035 691.725 10.365 ;
        RECT 691.395 8.675 691.725 9.005 ;
        RECT 691.395 7.315 691.725 7.645 ;
        RECT 691.395 5.955 691.725 6.285 ;
        RECT 691.395 4.595 691.725 4.925 ;
        RECT 691.395 3.235 691.725 3.565 ;
        RECT 691.395 1.875 691.725 2.205 ;
        RECT 691.395 0.515 691.725 0.845 ;
        RECT 691.4 -8.32 691.72 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 692.755 15.475 693.085 15.805 ;
        RECT 692.755 10.035 693.085 10.365 ;
        RECT 692.755 8.675 693.085 9.005 ;
        RECT 692.755 7.315 693.085 7.645 ;
        RECT 692.755 5.955 693.085 6.285 ;
        RECT 692.755 4.595 693.085 4.925 ;
        RECT 692.755 3.235 693.085 3.565 ;
        RECT 692.755 1.875 693.085 2.205 ;
        RECT 692.755 0.515 693.085 0.845 ;
        RECT 692.76 -8.32 693.08 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 694.115 15.475 694.445 15.805 ;
        RECT 694.115 10.035 694.445 10.365 ;
        RECT 694.115 8.675 694.445 9.005 ;
        RECT 694.115 7.315 694.445 7.645 ;
        RECT 694.115 5.955 694.445 6.285 ;
        RECT 694.115 4.595 694.445 4.925 ;
        RECT 694.115 3.235 694.445 3.565 ;
        RECT 694.115 1.875 694.445 2.205 ;
        RECT 694.115 0.515 694.445 0.845 ;
        RECT 694.12 -8.32 694.44 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 695.475 15.475 695.805 15.805 ;
        RECT 695.475 10.035 695.805 10.365 ;
        RECT 695.475 8.675 695.805 9.005 ;
        RECT 695.475 7.315 695.805 7.645 ;
        RECT 695.475 5.955 695.805 6.285 ;
        RECT 695.475 4.595 695.805 4.925 ;
        RECT 695.475 3.235 695.805 3.565 ;
        RECT 695.475 1.875 695.805 2.205 ;
        RECT 695.475 0.515 695.805 0.845 ;
        RECT 695.48 -8.32 695.8 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 696.835 15.475 697.165 15.805 ;
        RECT 696.835 10.035 697.165 10.365 ;
        RECT 696.835 8.675 697.165 9.005 ;
        RECT 696.835 7.315 697.165 7.645 ;
        RECT 696.835 5.955 697.165 6.285 ;
        RECT 696.835 4.595 697.165 4.925 ;
        RECT 696.835 3.235 697.165 3.565 ;
        RECT 696.835 1.875 697.165 2.205 ;
        RECT 696.835 0.515 697.165 0.845 ;
        RECT 696.84 -8.32 697.16 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 698.195 15.475 698.525 15.805 ;
        RECT 698.195 10.035 698.525 10.365 ;
        RECT 698.195 8.675 698.525 9.005 ;
        RECT 698.195 7.315 698.525 7.645 ;
        RECT 698.195 5.955 698.525 6.285 ;
        RECT 698.195 4.595 698.525 4.925 ;
        RECT 698.195 3.235 698.525 3.565 ;
        RECT 698.195 1.875 698.525 2.205 ;
        RECT 698.195 0.515 698.525 0.845 ;
        RECT 698.2 -8.32 698.52 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 699.555 15.475 699.885 15.805 ;
        RECT 699.555 11.395 699.885 11.725 ;
        RECT 699.555 10.035 699.885 10.365 ;
        RECT 699.555 8.675 699.885 9.005 ;
        RECT 699.555 7.315 699.885 7.645 ;
        RECT 699.555 5.955 699.885 6.285 ;
        RECT 699.555 4.595 699.885 4.925 ;
        RECT 699.555 3.235 699.885 3.565 ;
        RECT 699.555 1.875 699.885 2.205 ;
        RECT 699.555 0.515 699.885 0.845 ;
        RECT 699.56 -8.32 699.88 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 700.915 15.475 701.245 15.805 ;
        RECT 700.915 11.395 701.245 11.725 ;
        RECT 700.915 10.035 701.245 10.365 ;
        RECT 700.915 8.675 701.245 9.005 ;
        RECT 700.915 7.315 701.245 7.645 ;
        RECT 700.915 5.955 701.245 6.285 ;
        RECT 700.915 4.595 701.245 4.925 ;
        RECT 700.915 3.235 701.245 3.565 ;
        RECT 700.915 1.875 701.245 2.205 ;
        RECT 700.915 0.515 701.245 0.845 ;
        RECT 700.92 -8.32 701.24 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 702.275 15.475 702.605 15.805 ;
        RECT 702.275 11.395 702.605 11.725 ;
        RECT 702.275 10.035 702.605 10.365 ;
        RECT 702.275 8.675 702.605 9.005 ;
        RECT 702.275 7.315 702.605 7.645 ;
        RECT 702.275 5.955 702.605 6.285 ;
        RECT 702.275 4.595 702.605 4.925 ;
        RECT 702.275 3.235 702.605 3.565 ;
        RECT 702.275 1.875 702.605 2.205 ;
        RECT 702.275 0.515 702.605 0.845 ;
        RECT 702.28 -8.32 702.6 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 703.635 15.475 703.965 15.805 ;
        RECT 703.635 10.035 703.965 10.365 ;
        RECT 703.635 8.675 703.965 9.005 ;
        RECT 703.635 7.315 703.965 7.645 ;
        RECT 703.635 5.955 703.965 6.285 ;
        RECT 703.635 4.595 703.965 4.925 ;
        RECT 703.635 3.235 703.965 3.565 ;
        RECT 703.635 1.875 703.965 2.205 ;
        RECT 703.635 0.515 703.965 0.845 ;
        RECT 703.64 -8.32 703.96 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 704.995 15.475 705.325 15.805 ;
        RECT 704.995 10.035 705.325 10.365 ;
        RECT 704.995 8.675 705.325 9.005 ;
        RECT 704.995 7.315 705.325 7.645 ;
        RECT 704.995 5.955 705.325 6.285 ;
        RECT 704.995 4.595 705.325 4.925 ;
        RECT 704.995 3.235 705.325 3.565 ;
        RECT 704.995 1.875 705.325 2.205 ;
        RECT 704.995 0.515 705.325 0.845 ;
        RECT 705 -8.32 705.32 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 706.355 15.475 706.685 15.805 ;
        RECT 706.355 10.035 706.685 10.365 ;
        RECT 706.355 8.675 706.685 9.005 ;
        RECT 706.355 7.315 706.685 7.645 ;
        RECT 706.355 5.955 706.685 6.285 ;
        RECT 706.355 4.595 706.685 4.925 ;
        RECT 706.355 3.235 706.685 3.565 ;
        RECT 706.355 1.875 706.685 2.205 ;
        RECT 706.355 0.515 706.685 0.845 ;
        RECT 706.36 -8.32 706.68 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 707.715 15.475 708.045 15.805 ;
        RECT 707.715 10.035 708.045 10.365 ;
        RECT 707.715 8.675 708.045 9.005 ;
        RECT 707.715 7.315 708.045 7.645 ;
        RECT 707.715 5.955 708.045 6.285 ;
        RECT 707.715 4.595 708.045 4.925 ;
        RECT 707.715 3.235 708.045 3.565 ;
        RECT 707.715 1.875 708.045 2.205 ;
        RECT 707.715 0.515 708.045 0.845 ;
        RECT 707.72 -8.32 708.04 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 709.075 15.475 709.405 15.805 ;
        RECT 709.075 10.035 709.405 10.365 ;
        RECT 709.075 8.675 709.405 9.005 ;
        RECT 709.075 7.315 709.405 7.645 ;
        RECT 709.075 5.955 709.405 6.285 ;
        RECT 709.075 4.595 709.405 4.925 ;
        RECT 709.075 3.235 709.405 3.565 ;
        RECT 709.075 1.875 709.405 2.205 ;
        RECT 709.075 0.515 709.405 0.845 ;
        RECT 709.08 -8.32 709.4 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 710.435 15.475 710.765 15.805 ;
        RECT 710.435 10.035 710.765 10.365 ;
        RECT 710.435 8.675 710.765 9.005 ;
        RECT 710.435 7.315 710.765 7.645 ;
        RECT 710.435 5.955 710.765 6.285 ;
        RECT 710.435 4.595 710.765 4.925 ;
        RECT 710.435 3.235 710.765 3.565 ;
        RECT 710.435 1.875 710.765 2.205 ;
        RECT 710.435 0.515 710.765 0.845 ;
        RECT 710.44 -8.32 710.76 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 711.795 15.475 712.125 15.805 ;
        RECT 711.795 11.395 712.125 11.725 ;
        RECT 711.795 10.035 712.125 10.365 ;
        RECT 711.795 8.675 712.125 9.005 ;
        RECT 711.795 7.315 712.125 7.645 ;
        RECT 711.795 5.955 712.125 6.285 ;
        RECT 711.795 4.595 712.125 4.925 ;
        RECT 711.795 3.235 712.125 3.565 ;
        RECT 711.795 1.875 712.125 2.205 ;
        RECT 711.795 0.515 712.125 0.845 ;
        RECT 711.8 -8.32 712.12 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 713.155 15.475 713.485 15.805 ;
        RECT 713.155 11.395 713.485 11.725 ;
        RECT 713.155 10.035 713.485 10.365 ;
        RECT 713.155 8.675 713.485 9.005 ;
        RECT 713.155 7.315 713.485 7.645 ;
        RECT 713.155 5.955 713.485 6.285 ;
        RECT 713.155 4.595 713.485 4.925 ;
        RECT 713.155 3.235 713.485 3.565 ;
        RECT 713.155 1.875 713.485 2.205 ;
        RECT 713.155 0.515 713.485 0.845 ;
        RECT 713.16 -8.32 713.48 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 714.515 15.475 714.845 15.805 ;
        RECT 714.515 11.395 714.845 11.725 ;
        RECT 714.515 10.035 714.845 10.365 ;
        RECT 714.515 8.675 714.845 9.005 ;
        RECT 714.515 7.315 714.845 7.645 ;
        RECT 714.515 5.955 714.845 6.285 ;
        RECT 714.515 4.595 714.845 4.925 ;
        RECT 714.515 3.235 714.845 3.565 ;
        RECT 714.515 1.875 714.845 2.205 ;
        RECT 714.515 0.515 714.845 0.845 ;
        RECT 714.52 -8.32 714.84 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 715.875 15.475 716.205 15.805 ;
        RECT 715.875 10.035 716.205 10.365 ;
        RECT 715.875 8.675 716.205 9.005 ;
        RECT 715.875 7.315 716.205 7.645 ;
        RECT 715.875 5.955 716.205 6.285 ;
        RECT 715.875 4.595 716.205 4.925 ;
        RECT 715.875 3.235 716.205 3.565 ;
        RECT 715.875 1.875 716.205 2.205 ;
        RECT 715.875 0.515 716.205 0.845 ;
        RECT 715.88 -8.32 716.2 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 717.235 15.475 717.565 15.805 ;
        RECT 717.235 10.035 717.565 10.365 ;
        RECT 717.235 8.675 717.565 9.005 ;
        RECT 717.235 7.315 717.565 7.645 ;
        RECT 717.235 5.955 717.565 6.285 ;
        RECT 717.235 4.595 717.565 4.925 ;
        RECT 717.235 3.235 717.565 3.565 ;
        RECT 717.235 1.875 717.565 2.205 ;
        RECT 717.235 0.515 717.565 0.845 ;
        RECT 717.24 -8.32 717.56 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 718.595 15.475 718.925 15.805 ;
        RECT 718.595 10.035 718.925 10.365 ;
        RECT 718.595 8.675 718.925 9.005 ;
        RECT 718.595 7.315 718.925 7.645 ;
        RECT 718.595 5.955 718.925 6.285 ;
        RECT 718.595 4.595 718.925 4.925 ;
        RECT 718.595 3.235 718.925 3.565 ;
        RECT 718.595 1.875 718.925 2.205 ;
        RECT 718.595 0.515 718.925 0.845 ;
        RECT 718.6 -8.32 718.92 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 719.955 15.475 720.285 15.805 ;
        RECT 719.955 10.035 720.285 10.365 ;
        RECT 719.955 8.675 720.285 9.005 ;
        RECT 719.955 7.315 720.285 7.645 ;
        RECT 719.955 5.955 720.285 6.285 ;
        RECT 719.955 4.595 720.285 4.925 ;
        RECT 719.955 3.235 720.285 3.565 ;
        RECT 719.955 1.875 720.285 2.205 ;
        RECT 719.955 0.515 720.285 0.845 ;
        RECT 719.96 -8.32 720.28 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 721.315 15.475 721.645 15.805 ;
        RECT 721.315 10.035 721.645 10.365 ;
        RECT 721.315 8.675 721.645 9.005 ;
        RECT 721.315 7.315 721.645 7.645 ;
        RECT 721.315 5.955 721.645 6.285 ;
        RECT 721.315 4.595 721.645 4.925 ;
        RECT 721.315 3.235 721.645 3.565 ;
        RECT 721.315 1.875 721.645 2.205 ;
        RECT 721.315 0.515 721.645 0.845 ;
        RECT 721.32 -8.32 721.64 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 722.675 15.475 723.005 15.805 ;
        RECT 722.675 10.035 723.005 10.365 ;
        RECT 722.675 8.675 723.005 9.005 ;
        RECT 722.675 7.315 723.005 7.645 ;
        RECT 722.675 5.955 723.005 6.285 ;
        RECT 722.675 4.595 723.005 4.925 ;
        RECT 722.675 3.235 723.005 3.565 ;
        RECT 722.675 1.875 723.005 2.205 ;
        RECT 722.675 0.515 723.005 0.845 ;
        RECT 722.68 -8.32 723 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 724.035 15.475 724.365 15.805 ;
        RECT 724.035 11.395 724.365 11.725 ;
        RECT 724.035 10.035 724.365 10.365 ;
        RECT 724.035 8.675 724.365 9.005 ;
        RECT 724.035 7.315 724.365 7.645 ;
        RECT 724.035 5.955 724.365 6.285 ;
        RECT 724.035 4.595 724.365 4.925 ;
        RECT 724.035 3.235 724.365 3.565 ;
        RECT 724.035 1.875 724.365 2.205 ;
        RECT 724.035 0.515 724.365 0.845 ;
        RECT 724.04 -8.32 724.36 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 725.395 15.475 725.725 15.805 ;
        RECT 725.395 11.395 725.725 11.725 ;
        RECT 725.395 10.035 725.725 10.365 ;
        RECT 725.395 8.675 725.725 9.005 ;
        RECT 725.395 7.315 725.725 7.645 ;
        RECT 725.395 5.955 725.725 6.285 ;
        RECT 725.395 4.595 725.725 4.925 ;
        RECT 725.395 3.235 725.725 3.565 ;
        RECT 725.395 1.875 725.725 2.205 ;
        RECT 725.395 0.515 725.725 0.845 ;
        RECT 725.4 -8.32 725.72 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 726.755 15.475 727.085 15.805 ;
        RECT 726.755 11.395 727.085 11.725 ;
        RECT 726.755 10.035 727.085 10.365 ;
        RECT 726.755 8.675 727.085 9.005 ;
        RECT 726.755 7.315 727.085 7.645 ;
        RECT 726.755 5.955 727.085 6.285 ;
        RECT 726.755 4.595 727.085 4.925 ;
        RECT 726.755 3.235 727.085 3.565 ;
        RECT 726.755 1.875 727.085 2.205 ;
        RECT 726.755 0.515 727.085 0.845 ;
        RECT 726.76 -8.32 727.08 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 728.115 15.475 728.445 15.805 ;
        RECT 728.115 10.035 728.445 10.365 ;
        RECT 728.115 8.675 728.445 9.005 ;
        RECT 728.115 7.315 728.445 7.645 ;
        RECT 728.115 5.955 728.445 6.285 ;
        RECT 728.115 4.595 728.445 4.925 ;
        RECT 728.115 3.235 728.445 3.565 ;
        RECT 728.115 1.875 728.445 2.205 ;
        RECT 728.115 0.515 728.445 0.845 ;
        RECT 728.12 -8.32 728.44 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 729.475 15.475 729.805 15.805 ;
        RECT 729.475 10.035 729.805 10.365 ;
        RECT 729.475 8.675 729.805 9.005 ;
        RECT 729.475 7.315 729.805 7.645 ;
        RECT 729.475 5.955 729.805 6.285 ;
        RECT 729.475 4.595 729.805 4.925 ;
        RECT 729.475 3.235 729.805 3.565 ;
        RECT 729.475 1.875 729.805 2.205 ;
        RECT 729.475 0.515 729.805 0.845 ;
        RECT 729.48 -8.32 729.8 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 730.835 15.475 731.165 15.805 ;
        RECT 730.835 10.035 731.165 10.365 ;
        RECT 730.835 8.675 731.165 9.005 ;
        RECT 730.835 7.315 731.165 7.645 ;
        RECT 730.835 5.955 731.165 6.285 ;
        RECT 730.835 4.595 731.165 4.925 ;
        RECT 730.835 3.235 731.165 3.565 ;
        RECT 730.835 1.875 731.165 2.205 ;
        RECT 730.835 0.515 731.165 0.845 ;
        RECT 730.84 -8.32 731.16 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 732.195 15.475 732.525 15.805 ;
        RECT 732.195 10.035 732.525 10.365 ;
        RECT 732.195 8.675 732.525 9.005 ;
        RECT 732.195 7.315 732.525 7.645 ;
        RECT 732.195 5.955 732.525 6.285 ;
        RECT 732.195 4.595 732.525 4.925 ;
        RECT 732.195 3.235 732.525 3.565 ;
        RECT 732.195 1.875 732.525 2.205 ;
        RECT 732.195 0.515 732.525 0.845 ;
        RECT 732.2 -8.32 732.52 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 733.555 15.475 733.885 15.805 ;
        RECT 733.555 10.035 733.885 10.365 ;
        RECT 733.555 8.675 733.885 9.005 ;
        RECT 733.555 7.315 733.885 7.645 ;
        RECT 733.555 5.955 733.885 6.285 ;
        RECT 733.555 4.595 733.885 4.925 ;
        RECT 733.555 3.235 733.885 3.565 ;
        RECT 733.555 1.875 733.885 2.205 ;
        RECT 733.555 0.515 733.885 0.845 ;
        RECT 733.56 -8.32 733.88 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 734.915 15.475 735.245 15.805 ;
        RECT 734.915 11.395 735.245 11.725 ;
        RECT 734.915 10.035 735.245 10.365 ;
        RECT 734.915 8.675 735.245 9.005 ;
        RECT 734.915 7.315 735.245 7.645 ;
        RECT 734.915 5.955 735.245 6.285 ;
        RECT 734.915 4.595 735.245 4.925 ;
        RECT 734.915 3.235 735.245 3.565 ;
        RECT 734.915 1.875 735.245 2.205 ;
        RECT 734.915 0.515 735.245 0.845 ;
        RECT 734.92 -8.32 735.24 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 736.275 15.475 736.605 15.805 ;
        RECT 736.275 11.395 736.605 11.725 ;
        RECT 736.275 10.035 736.605 10.365 ;
        RECT 736.275 8.675 736.605 9.005 ;
        RECT 736.275 7.315 736.605 7.645 ;
        RECT 736.275 5.955 736.605 6.285 ;
        RECT 736.275 4.595 736.605 4.925 ;
        RECT 736.275 3.235 736.605 3.565 ;
        RECT 736.275 1.875 736.605 2.205 ;
        RECT 736.275 0.515 736.605 0.845 ;
        RECT 736.28 -8.32 736.6 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 737.635 15.475 737.965 15.805 ;
        RECT 737.635 11.395 737.965 11.725 ;
        RECT 737.635 10.035 737.965 10.365 ;
        RECT 737.635 8.675 737.965 9.005 ;
        RECT 737.635 7.315 737.965 7.645 ;
        RECT 737.635 5.955 737.965 6.285 ;
        RECT 737.635 4.595 737.965 4.925 ;
        RECT 737.635 3.235 737.965 3.565 ;
        RECT 737.635 1.875 737.965 2.205 ;
        RECT 737.635 0.515 737.965 0.845 ;
        RECT 737.64 -8.32 737.96 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 738.995 15.475 739.325 15.805 ;
        RECT 738.995 10.035 739.325 10.365 ;
        RECT 738.995 8.675 739.325 9.005 ;
        RECT 738.995 7.315 739.325 7.645 ;
        RECT 738.995 5.955 739.325 6.285 ;
        RECT 738.995 4.595 739.325 4.925 ;
        RECT 738.995 3.235 739.325 3.565 ;
        RECT 738.995 1.875 739.325 2.205 ;
        RECT 738.995 0.515 739.325 0.845 ;
        RECT 739 -8.32 739.32 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 740.355 15.475 740.685 15.805 ;
        RECT 740.355 10.035 740.685 10.365 ;
        RECT 740.355 8.675 740.685 9.005 ;
        RECT 740.355 7.315 740.685 7.645 ;
        RECT 740.355 5.955 740.685 6.285 ;
        RECT 740.355 4.595 740.685 4.925 ;
        RECT 740.355 3.235 740.685 3.565 ;
        RECT 740.355 1.875 740.685 2.205 ;
        RECT 740.355 0.515 740.685 0.845 ;
        RECT 740.36 -8.32 740.68 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 741.715 15.475 742.045 15.805 ;
        RECT 741.715 10.035 742.045 10.365 ;
        RECT 741.715 8.675 742.045 9.005 ;
        RECT 741.715 7.315 742.045 7.645 ;
        RECT 741.715 5.955 742.045 6.285 ;
        RECT 741.715 4.595 742.045 4.925 ;
        RECT 741.715 3.235 742.045 3.565 ;
        RECT 741.715 1.875 742.045 2.205 ;
        RECT 741.715 0.515 742.045 0.845 ;
        RECT 741.72 -8.32 742.04 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 743.075 15.475 743.405 15.805 ;
        RECT 743.075 10.035 743.405 10.365 ;
        RECT 743.075 8.675 743.405 9.005 ;
        RECT 743.075 7.315 743.405 7.645 ;
        RECT 743.075 5.955 743.405 6.285 ;
        RECT 743.075 4.595 743.405 4.925 ;
        RECT 743.075 3.235 743.405 3.565 ;
        RECT 743.075 1.875 743.405 2.205 ;
        RECT 743.075 0.515 743.405 0.845 ;
        RECT 743.08 -8.32 743.4 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 744.435 15.475 744.765 15.805 ;
        RECT 744.435 10.035 744.765 10.365 ;
        RECT 744.435 8.675 744.765 9.005 ;
        RECT 744.435 7.315 744.765 7.645 ;
        RECT 744.435 5.955 744.765 6.285 ;
        RECT 744.435 4.595 744.765 4.925 ;
        RECT 744.435 3.235 744.765 3.565 ;
        RECT 744.435 1.875 744.765 2.205 ;
        RECT 744.435 0.515 744.765 0.845 ;
        RECT 744.44 -8.32 744.76 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 745.795 15.475 746.125 15.805 ;
        RECT 745.795 10.035 746.125 10.365 ;
        RECT 745.795 8.675 746.125 9.005 ;
        RECT 745.795 7.315 746.125 7.645 ;
        RECT 745.795 5.955 746.125 6.285 ;
        RECT 745.795 4.595 746.125 4.925 ;
        RECT 745.795 3.235 746.125 3.565 ;
        RECT 745.795 1.875 746.125 2.205 ;
        RECT 745.795 0.515 746.125 0.845 ;
        RECT 745.8 -8.32 746.12 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 747.155 15.475 747.485 15.805 ;
        RECT 747.155 11.395 747.485 11.725 ;
        RECT 747.155 10.035 747.485 10.365 ;
        RECT 747.155 8.675 747.485 9.005 ;
        RECT 747.155 7.315 747.485 7.645 ;
        RECT 747.155 5.955 747.485 6.285 ;
        RECT 747.155 4.595 747.485 4.925 ;
        RECT 747.155 3.235 747.485 3.565 ;
        RECT 747.155 1.875 747.485 2.205 ;
        RECT 747.155 0.515 747.485 0.845 ;
        RECT 747.16 -8.32 747.48 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 748.515 15.475 748.845 15.805 ;
        RECT 748.515 11.395 748.845 11.725 ;
        RECT 748.515 10.035 748.845 10.365 ;
        RECT 748.515 8.675 748.845 9.005 ;
        RECT 748.515 7.315 748.845 7.645 ;
        RECT 748.515 5.955 748.845 6.285 ;
        RECT 748.515 4.595 748.845 4.925 ;
        RECT 748.515 3.235 748.845 3.565 ;
        RECT 748.515 1.875 748.845 2.205 ;
        RECT 748.515 0.515 748.845 0.845 ;
        RECT 748.52 -8.32 748.84 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 749.875 15.475 750.205 15.805 ;
        RECT 749.875 11.395 750.205 11.725 ;
        RECT 749.875 10.035 750.205 10.365 ;
        RECT 749.875 8.675 750.205 9.005 ;
        RECT 749.875 7.315 750.205 7.645 ;
        RECT 749.875 5.955 750.205 6.285 ;
        RECT 749.875 4.595 750.205 4.925 ;
        RECT 749.875 3.235 750.205 3.565 ;
        RECT 749.875 1.875 750.205 2.205 ;
        RECT 749.875 0.515 750.205 0.845 ;
        RECT 749.88 -8.32 750.2 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 751.235 15.475 751.565 15.805 ;
        RECT 751.235 10.035 751.565 10.365 ;
        RECT 751.235 8.675 751.565 9.005 ;
        RECT 751.235 7.315 751.565 7.645 ;
        RECT 751.235 5.955 751.565 6.285 ;
        RECT 751.235 4.595 751.565 4.925 ;
        RECT 751.235 3.235 751.565 3.565 ;
        RECT 751.235 1.875 751.565 2.205 ;
        RECT 751.235 0.515 751.565 0.845 ;
        RECT 751.24 -8.32 751.56 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 752.595 15.475 752.925 15.805 ;
        RECT 752.595 10.035 752.925 10.365 ;
        RECT 752.595 8.675 752.925 9.005 ;
        RECT 752.595 7.315 752.925 7.645 ;
        RECT 752.595 5.955 752.925 6.285 ;
        RECT 752.595 4.595 752.925 4.925 ;
        RECT 752.595 3.235 752.925 3.565 ;
        RECT 752.595 1.875 752.925 2.205 ;
        RECT 752.595 0.515 752.925 0.845 ;
        RECT 752.6 -8.32 752.92 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 753.955 15.475 754.285 15.805 ;
        RECT 753.955 10.035 754.285 10.365 ;
        RECT 753.955 8.675 754.285 9.005 ;
        RECT 753.955 7.315 754.285 7.645 ;
        RECT 753.955 5.955 754.285 6.285 ;
        RECT 753.955 4.595 754.285 4.925 ;
        RECT 753.955 3.235 754.285 3.565 ;
        RECT 753.955 1.875 754.285 2.205 ;
        RECT 753.955 0.515 754.285 0.845 ;
        RECT 753.96 -8.32 754.28 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 755.315 15.475 755.645 15.805 ;
        RECT 755.315 10.035 755.645 10.365 ;
        RECT 755.315 8.675 755.645 9.005 ;
        RECT 755.315 7.315 755.645 7.645 ;
        RECT 755.315 5.955 755.645 6.285 ;
        RECT 755.315 4.595 755.645 4.925 ;
        RECT 755.315 3.235 755.645 3.565 ;
        RECT 755.315 1.875 755.645 2.205 ;
        RECT 755.315 0.515 755.645 0.845 ;
        RECT 755.32 -8.32 755.64 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 756.675 15.475 757.005 15.805 ;
        RECT 756.675 10.035 757.005 10.365 ;
        RECT 756.675 8.675 757.005 9.005 ;
        RECT 756.675 7.315 757.005 7.645 ;
        RECT 756.675 5.955 757.005 6.285 ;
        RECT 756.675 4.595 757.005 4.925 ;
        RECT 756.675 3.235 757.005 3.565 ;
        RECT 756.675 1.875 757.005 2.205 ;
        RECT 756.675 0.515 757.005 0.845 ;
        RECT 756.68 -8.32 757 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 758.035 15.475 758.365 15.805 ;
        RECT 758.035 10.035 758.365 10.365 ;
        RECT 758.035 8.675 758.365 9.005 ;
        RECT 758.035 7.315 758.365 7.645 ;
        RECT 758.035 5.955 758.365 6.285 ;
        RECT 758.035 4.595 758.365 4.925 ;
        RECT 758.035 3.235 758.365 3.565 ;
        RECT 758.035 1.875 758.365 2.205 ;
        RECT 758.035 0.515 758.365 0.845 ;
        RECT 758.04 -8.32 758.36 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 759.395 15.475 759.725 15.805 ;
        RECT 759.395 11.395 759.725 11.725 ;
        RECT 759.395 10.035 759.725 10.365 ;
        RECT 759.395 8.675 759.725 9.005 ;
        RECT 759.395 7.315 759.725 7.645 ;
        RECT 759.395 5.955 759.725 6.285 ;
        RECT 759.395 4.595 759.725 4.925 ;
        RECT 759.395 3.235 759.725 3.565 ;
        RECT 759.395 1.875 759.725 2.205 ;
        RECT 759.395 0.515 759.725 0.845 ;
        RECT 759.4 -8.32 759.72 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 760.755 15.475 761.085 15.805 ;
        RECT 760.755 11.395 761.085 11.725 ;
        RECT 760.755 10.035 761.085 10.365 ;
        RECT 760.755 8.675 761.085 9.005 ;
        RECT 760.755 7.315 761.085 7.645 ;
        RECT 760.755 5.955 761.085 6.285 ;
        RECT 760.755 4.595 761.085 4.925 ;
        RECT 760.755 3.235 761.085 3.565 ;
        RECT 760.755 1.875 761.085 2.205 ;
        RECT 760.755 0.515 761.085 0.845 ;
        RECT 760.76 -8.32 761.08 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 762.115 15.475 762.445 15.805 ;
        RECT 762.115 11.395 762.445 11.725 ;
        RECT 762.115 10.035 762.445 10.365 ;
        RECT 762.115 8.675 762.445 9.005 ;
        RECT 762.115 7.315 762.445 7.645 ;
        RECT 762.115 5.955 762.445 6.285 ;
        RECT 762.115 4.595 762.445 4.925 ;
        RECT 762.115 3.235 762.445 3.565 ;
        RECT 762.115 1.875 762.445 2.205 ;
        RECT 762.115 0.515 762.445 0.845 ;
        RECT 762.12 -8.32 762.44 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 763.475 15.475 763.805 15.805 ;
        RECT 763.475 11.395 763.805 11.725 ;
        RECT 763.475 10.035 763.805 10.365 ;
        RECT 763.475 8.675 763.805 9.005 ;
        RECT 763.475 7.315 763.805 7.645 ;
        RECT 763.475 5.955 763.805 6.285 ;
        RECT 763.475 4.595 763.805 4.925 ;
        RECT 763.475 3.235 763.805 3.565 ;
        RECT 763.475 1.875 763.805 2.205 ;
        RECT 763.475 0.515 763.805 0.845 ;
        RECT 763.48 -8.32 763.8 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 764.835 15.475 765.165 15.805 ;
        RECT 764.835 12.755 765.165 13.085 ;
        RECT 764.835 11.395 765.165 11.725 ;
        RECT 764.835 10.035 765.165 10.365 ;
        RECT 764.835 8.675 765.165 9.005 ;
        RECT 764.835 7.315 765.165 7.645 ;
        RECT 764.835 5.955 765.165 6.285 ;
        RECT 764.835 4.595 765.165 4.925 ;
        RECT 764.835 3.235 765.165 3.565 ;
        RECT 764.835 1.875 765.165 2.205 ;
        RECT 764.835 0.515 765.165 0.845 ;
        RECT 764.84 -8.32 765.16 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 766.195 15.475 766.525 15.805 ;
        RECT 766.195 12.755 766.525 13.085 ;
        RECT 766.195 11.395 766.525 11.725 ;
        RECT 766.195 10.035 766.525 10.365 ;
        RECT 766.195 8.675 766.525 9.005 ;
        RECT 766.195 7.315 766.525 7.645 ;
        RECT 766.195 5.955 766.525 6.285 ;
        RECT 766.195 4.595 766.525 4.925 ;
        RECT 766.195 3.235 766.525 3.565 ;
        RECT 766.195 1.875 766.525 2.205 ;
        RECT 766.195 0.515 766.525 0.845 ;
        RECT 766.2 -8.32 766.52 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 767.555 15.475 767.885 15.805 ;
        RECT 767.555 14.115 767.885 14.445 ;
        RECT 767.555 12.755 767.885 13.085 ;
        RECT 767.555 11.395 767.885 11.725 ;
        RECT 767.555 10.035 767.885 10.365 ;
        RECT 767.555 8.675 767.885 9.005 ;
        RECT 767.555 7.315 767.885 7.645 ;
        RECT 767.555 5.955 767.885 6.285 ;
        RECT 767.555 4.595 767.885 4.925 ;
        RECT 767.555 3.235 767.885 3.565 ;
        RECT 767.555 1.875 767.885 2.205 ;
        RECT 767.555 0.515 767.885 0.845 ;
        RECT 767.56 -8.32 767.88 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 768.915 15.475 769.245 15.805 ;
        RECT 768.915 14.115 769.245 14.445 ;
        RECT 768.915 12.755 769.245 13.085 ;
        RECT 768.915 11.395 769.245 11.725 ;
        RECT 768.915 10.035 769.245 10.365 ;
        RECT 768.915 8.675 769.245 9.005 ;
        RECT 768.915 7.315 769.245 7.645 ;
        RECT 768.915 5.955 769.245 6.285 ;
        RECT 768.915 4.595 769.245 4.925 ;
        RECT 768.915 3.235 769.245 3.565 ;
        RECT 768.915 1.875 769.245 2.205 ;
        RECT 768.915 0.515 769.245 0.845 ;
        RECT 768.92 -8.32 769.24 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 509.155 15.475 509.485 15.805 ;
        RECT 509.155 11.395 509.485 11.725 ;
        RECT 509.155 10.035 509.485 10.365 ;
        RECT 509.155 8.675 509.485 9.005 ;
        RECT 509.155 7.315 509.485 7.645 ;
        RECT 509.155 5.955 509.485 6.285 ;
        RECT 509.155 4.595 509.485 4.925 ;
        RECT 509.155 3.235 509.485 3.565 ;
        RECT 509.155 1.875 509.485 2.205 ;
        RECT 509.155 0.515 509.485 0.845 ;
        RECT 509.16 -8.32 509.48 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 510.515 15.475 510.845 15.805 ;
        RECT 510.515 11.395 510.845 11.725 ;
        RECT 510.515 10.035 510.845 10.365 ;
        RECT 510.515 8.675 510.845 9.005 ;
        RECT 510.515 7.315 510.845 7.645 ;
        RECT 510.515 5.955 510.845 6.285 ;
        RECT 510.515 4.595 510.845 4.925 ;
        RECT 510.515 3.235 510.845 3.565 ;
        RECT 510.515 1.875 510.845 2.205 ;
        RECT 510.515 0.515 510.845 0.845 ;
        RECT 510.52 -8.32 510.84 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 511.875 15.475 512.205 15.805 ;
        RECT 511.875 10.035 512.205 10.365 ;
        RECT 511.875 8.675 512.205 9.005 ;
        RECT 511.875 7.315 512.205 7.645 ;
        RECT 511.875 5.955 512.205 6.285 ;
        RECT 511.875 4.595 512.205 4.925 ;
        RECT 511.875 3.235 512.205 3.565 ;
        RECT 511.875 1.875 512.205 2.205 ;
        RECT 511.875 0.515 512.205 0.845 ;
        RECT 511.88 -8.32 512.2 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 513.235 15.475 513.565 15.805 ;
        RECT 513.235 10.035 513.565 10.365 ;
        RECT 513.235 8.675 513.565 9.005 ;
        RECT 513.235 7.315 513.565 7.645 ;
        RECT 513.235 5.955 513.565 6.285 ;
        RECT 513.235 4.595 513.565 4.925 ;
        RECT 513.235 3.235 513.565 3.565 ;
        RECT 513.235 1.875 513.565 2.205 ;
        RECT 513.235 0.515 513.565 0.845 ;
        RECT 513.24 -8.32 513.56 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 514.595 15.475 514.925 15.805 ;
        RECT 514.595 10.035 514.925 10.365 ;
        RECT 514.595 8.675 514.925 9.005 ;
        RECT 514.595 7.315 514.925 7.645 ;
        RECT 514.595 5.955 514.925 6.285 ;
        RECT 514.595 4.595 514.925 4.925 ;
        RECT 514.595 3.235 514.925 3.565 ;
        RECT 514.595 1.875 514.925 2.205 ;
        RECT 514.595 0.515 514.925 0.845 ;
        RECT 514.6 -8.32 514.92 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 515.955 15.475 516.285 15.805 ;
        RECT 515.955 10.035 516.285 10.365 ;
        RECT 515.955 8.675 516.285 9.005 ;
        RECT 515.955 7.315 516.285 7.645 ;
        RECT 515.955 5.955 516.285 6.285 ;
        RECT 515.955 4.595 516.285 4.925 ;
        RECT 515.955 3.235 516.285 3.565 ;
        RECT 515.955 1.875 516.285 2.205 ;
        RECT 515.955 0.515 516.285 0.845 ;
        RECT 515.96 -8.32 516.28 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 517.315 15.475 517.645 15.805 ;
        RECT 517.315 10.035 517.645 10.365 ;
        RECT 517.315 8.675 517.645 9.005 ;
        RECT 517.315 7.315 517.645 7.645 ;
        RECT 517.315 5.955 517.645 6.285 ;
        RECT 517.315 4.595 517.645 4.925 ;
        RECT 517.315 3.235 517.645 3.565 ;
        RECT 517.315 1.875 517.645 2.205 ;
        RECT 517.315 0.515 517.645 0.845 ;
        RECT 517.32 -8.32 517.64 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 518.675 15.475 519.005 15.805 ;
        RECT 518.675 10.035 519.005 10.365 ;
        RECT 518.675 8.675 519.005 9.005 ;
        RECT 518.675 7.315 519.005 7.645 ;
        RECT 518.675 5.955 519.005 6.285 ;
        RECT 518.675 4.595 519.005 4.925 ;
        RECT 518.675 3.235 519.005 3.565 ;
        RECT 518.675 1.875 519.005 2.205 ;
        RECT 518.675 0.515 519.005 0.845 ;
        RECT 518.68 -8.32 519 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 520.035 15.475 520.365 15.805 ;
        RECT 520.035 11.395 520.365 11.725 ;
        RECT 520.035 10.035 520.365 10.365 ;
        RECT 520.035 8.675 520.365 9.005 ;
        RECT 520.035 7.315 520.365 7.645 ;
        RECT 520.035 5.955 520.365 6.285 ;
        RECT 520.035 4.595 520.365 4.925 ;
        RECT 520.035 3.235 520.365 3.565 ;
        RECT 520.035 1.875 520.365 2.205 ;
        RECT 520.035 0.515 520.365 0.845 ;
        RECT 520.04 -8.32 520.36 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 521.395 15.475 521.725 15.805 ;
        RECT 521.395 11.395 521.725 11.725 ;
        RECT 521.395 10.035 521.725 10.365 ;
        RECT 521.395 8.675 521.725 9.005 ;
        RECT 521.395 7.315 521.725 7.645 ;
        RECT 521.395 5.955 521.725 6.285 ;
        RECT 521.395 4.595 521.725 4.925 ;
        RECT 521.395 3.235 521.725 3.565 ;
        RECT 521.395 1.875 521.725 2.205 ;
        RECT 521.395 0.515 521.725 0.845 ;
        RECT 521.4 -8.32 521.72 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 522.755 15.475 523.085 15.805 ;
        RECT 522.755 11.395 523.085 11.725 ;
        RECT 522.755 10.035 523.085 10.365 ;
        RECT 522.755 8.675 523.085 9.005 ;
        RECT 522.755 7.315 523.085 7.645 ;
        RECT 522.755 5.955 523.085 6.285 ;
        RECT 522.755 4.595 523.085 4.925 ;
        RECT 522.755 3.235 523.085 3.565 ;
        RECT 522.755 1.875 523.085 2.205 ;
        RECT 522.755 0.515 523.085 0.845 ;
        RECT 522.76 -8.32 523.08 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 524.115 15.475 524.445 15.805 ;
        RECT 524.115 10.035 524.445 10.365 ;
        RECT 524.115 8.675 524.445 9.005 ;
        RECT 524.115 7.315 524.445 7.645 ;
        RECT 524.115 5.955 524.445 6.285 ;
        RECT 524.115 4.595 524.445 4.925 ;
        RECT 524.115 3.235 524.445 3.565 ;
        RECT 524.115 1.875 524.445 2.205 ;
        RECT 524.115 0.515 524.445 0.845 ;
        RECT 524.12 -8.32 524.44 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 525.475 15.475 525.805 15.805 ;
        RECT 525.475 10.035 525.805 10.365 ;
        RECT 525.475 8.675 525.805 9.005 ;
        RECT 525.475 7.315 525.805 7.645 ;
        RECT 525.475 5.955 525.805 6.285 ;
        RECT 525.475 4.595 525.805 4.925 ;
        RECT 525.475 3.235 525.805 3.565 ;
        RECT 525.475 1.875 525.805 2.205 ;
        RECT 525.475 0.515 525.805 0.845 ;
        RECT 525.48 -8.32 525.8 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 526.835 15.475 527.165 15.805 ;
        RECT 526.835 10.035 527.165 10.365 ;
        RECT 526.835 8.675 527.165 9.005 ;
        RECT 526.835 7.315 527.165 7.645 ;
        RECT 526.835 5.955 527.165 6.285 ;
        RECT 526.835 4.595 527.165 4.925 ;
        RECT 526.835 3.235 527.165 3.565 ;
        RECT 526.835 1.875 527.165 2.205 ;
        RECT 526.835 0.515 527.165 0.845 ;
        RECT 526.84 -8.32 527.16 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 528.195 15.475 528.525 15.805 ;
        RECT 528.195 10.035 528.525 10.365 ;
        RECT 528.195 8.675 528.525 9.005 ;
        RECT 528.195 7.315 528.525 7.645 ;
        RECT 528.195 5.955 528.525 6.285 ;
        RECT 528.195 4.595 528.525 4.925 ;
        RECT 528.195 3.235 528.525 3.565 ;
        RECT 528.195 1.875 528.525 2.205 ;
        RECT 528.195 0.515 528.525 0.845 ;
        RECT 528.2 -8.32 528.52 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 529.555 15.475 529.885 15.805 ;
        RECT 529.555 10.035 529.885 10.365 ;
        RECT 529.555 8.675 529.885 9.005 ;
        RECT 529.555 7.315 529.885 7.645 ;
        RECT 529.555 5.955 529.885 6.285 ;
        RECT 529.555 4.595 529.885 4.925 ;
        RECT 529.555 3.235 529.885 3.565 ;
        RECT 529.555 1.875 529.885 2.205 ;
        RECT 529.555 0.515 529.885 0.845 ;
        RECT 529.56 -8.32 529.88 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 530.915 15.475 531.245 15.805 ;
        RECT 530.915 11.395 531.245 11.725 ;
        RECT 530.915 10.035 531.245 10.365 ;
        RECT 530.915 8.675 531.245 9.005 ;
        RECT 530.915 7.315 531.245 7.645 ;
        RECT 530.915 5.955 531.245 6.285 ;
        RECT 530.915 4.595 531.245 4.925 ;
        RECT 530.915 3.235 531.245 3.565 ;
        RECT 530.915 1.875 531.245 2.205 ;
        RECT 530.915 0.515 531.245 0.845 ;
        RECT 530.92 -8.32 531.24 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 532.275 15.475 532.605 15.805 ;
        RECT 532.275 11.395 532.605 11.725 ;
        RECT 532.275 10.035 532.605 10.365 ;
        RECT 532.275 8.675 532.605 9.005 ;
        RECT 532.275 7.315 532.605 7.645 ;
        RECT 532.275 5.955 532.605 6.285 ;
        RECT 532.275 4.595 532.605 4.925 ;
        RECT 532.275 3.235 532.605 3.565 ;
        RECT 532.275 1.875 532.605 2.205 ;
        RECT 532.275 0.515 532.605 0.845 ;
        RECT 532.28 -8.32 532.6 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 533.635 15.475 533.965 15.805 ;
        RECT 533.635 11.395 533.965 11.725 ;
        RECT 533.635 10.035 533.965 10.365 ;
        RECT 533.635 8.675 533.965 9.005 ;
        RECT 533.635 7.315 533.965 7.645 ;
        RECT 533.635 5.955 533.965 6.285 ;
        RECT 533.635 4.595 533.965 4.925 ;
        RECT 533.635 3.235 533.965 3.565 ;
        RECT 533.635 1.875 533.965 2.205 ;
        RECT 533.635 0.515 533.965 0.845 ;
        RECT 533.64 -8.32 533.96 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 534.995 15.475 535.325 15.805 ;
        RECT 534.995 10.035 535.325 10.365 ;
        RECT 534.995 8.675 535.325 9.005 ;
        RECT 534.995 7.315 535.325 7.645 ;
        RECT 534.995 5.955 535.325 6.285 ;
        RECT 534.995 4.595 535.325 4.925 ;
        RECT 534.995 3.235 535.325 3.565 ;
        RECT 534.995 1.875 535.325 2.205 ;
        RECT 534.995 0.515 535.325 0.845 ;
        RECT 535 -8.32 535.32 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 536.355 15.475 536.685 15.805 ;
        RECT 536.355 10.035 536.685 10.365 ;
        RECT 536.355 8.675 536.685 9.005 ;
        RECT 536.355 7.315 536.685 7.645 ;
        RECT 536.355 5.955 536.685 6.285 ;
        RECT 536.355 4.595 536.685 4.925 ;
        RECT 536.355 3.235 536.685 3.565 ;
        RECT 536.355 1.875 536.685 2.205 ;
        RECT 536.355 0.515 536.685 0.845 ;
        RECT 536.36 -8.32 536.68 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 537.715 15.475 538.045 15.805 ;
        RECT 537.715 10.035 538.045 10.365 ;
        RECT 537.715 8.675 538.045 9.005 ;
        RECT 537.715 7.315 538.045 7.645 ;
        RECT 537.715 5.955 538.045 6.285 ;
        RECT 537.715 4.595 538.045 4.925 ;
        RECT 537.715 3.235 538.045 3.565 ;
        RECT 537.715 1.875 538.045 2.205 ;
        RECT 537.715 0.515 538.045 0.845 ;
        RECT 537.72 -8.32 538.04 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 539.075 15.475 539.405 15.805 ;
        RECT 539.075 10.035 539.405 10.365 ;
        RECT 539.075 8.675 539.405 9.005 ;
        RECT 539.075 7.315 539.405 7.645 ;
        RECT 539.075 5.955 539.405 6.285 ;
        RECT 539.075 4.595 539.405 4.925 ;
        RECT 539.075 3.235 539.405 3.565 ;
        RECT 539.075 1.875 539.405 2.205 ;
        RECT 539.075 0.515 539.405 0.845 ;
        RECT 539.08 -8.32 539.4 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 540.435 15.475 540.765 15.805 ;
        RECT 540.435 10.035 540.765 10.365 ;
        RECT 540.435 8.675 540.765 9.005 ;
        RECT 540.435 7.315 540.765 7.645 ;
        RECT 540.435 5.955 540.765 6.285 ;
        RECT 540.435 4.595 540.765 4.925 ;
        RECT 540.435 3.235 540.765 3.565 ;
        RECT 540.435 1.875 540.765 2.205 ;
        RECT 540.435 0.515 540.765 0.845 ;
        RECT 540.44 -8.32 540.76 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 541.795 15.475 542.125 15.805 ;
        RECT 541.795 10.035 542.125 10.365 ;
        RECT 541.795 8.675 542.125 9.005 ;
        RECT 541.795 7.315 542.125 7.645 ;
        RECT 541.795 5.955 542.125 6.285 ;
        RECT 541.795 4.595 542.125 4.925 ;
        RECT 541.795 3.235 542.125 3.565 ;
        RECT 541.795 1.875 542.125 2.205 ;
        RECT 541.795 0.515 542.125 0.845 ;
        RECT 541.8 -8.32 542.12 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 543.155 15.475 543.485 15.805 ;
        RECT 543.155 11.395 543.485 11.725 ;
        RECT 543.155 10.035 543.485 10.365 ;
        RECT 543.155 8.675 543.485 9.005 ;
        RECT 543.155 7.315 543.485 7.645 ;
        RECT 543.155 5.955 543.485 6.285 ;
        RECT 543.155 4.595 543.485 4.925 ;
        RECT 543.155 3.235 543.485 3.565 ;
        RECT 543.155 1.875 543.485 2.205 ;
        RECT 543.155 0.515 543.485 0.845 ;
        RECT 543.16 -8.32 543.48 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 544.515 15.475 544.845 15.805 ;
        RECT 544.515 11.395 544.845 11.725 ;
        RECT 544.515 10.035 544.845 10.365 ;
        RECT 544.515 8.675 544.845 9.005 ;
        RECT 544.515 7.315 544.845 7.645 ;
        RECT 544.515 5.955 544.845 6.285 ;
        RECT 544.515 4.595 544.845 4.925 ;
        RECT 544.515 3.235 544.845 3.565 ;
        RECT 544.515 1.875 544.845 2.205 ;
        RECT 544.515 0.515 544.845 0.845 ;
        RECT 544.52 -8.32 544.84 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 545.875 15.475 546.205 15.805 ;
        RECT 545.875 11.395 546.205 11.725 ;
        RECT 545.875 10.035 546.205 10.365 ;
        RECT 545.875 8.675 546.205 9.005 ;
        RECT 545.875 7.315 546.205 7.645 ;
        RECT 545.875 5.955 546.205 6.285 ;
        RECT 545.875 4.595 546.205 4.925 ;
        RECT 545.875 3.235 546.205 3.565 ;
        RECT 545.875 1.875 546.205 2.205 ;
        RECT 545.875 0.515 546.205 0.845 ;
        RECT 545.88 -8.32 546.2 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 547.235 15.475 547.565 15.805 ;
        RECT 547.235 10.035 547.565 10.365 ;
        RECT 547.235 8.675 547.565 9.005 ;
        RECT 547.235 7.315 547.565 7.645 ;
        RECT 547.235 5.955 547.565 6.285 ;
        RECT 547.235 4.595 547.565 4.925 ;
        RECT 547.235 3.235 547.565 3.565 ;
        RECT 547.235 1.875 547.565 2.205 ;
        RECT 547.235 0.515 547.565 0.845 ;
        RECT 547.24 -8.32 547.56 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 548.595 15.475 548.925 15.805 ;
        RECT 548.595 10.035 548.925 10.365 ;
        RECT 548.595 8.675 548.925 9.005 ;
        RECT 548.595 7.315 548.925 7.645 ;
        RECT 548.595 5.955 548.925 6.285 ;
        RECT 548.595 4.595 548.925 4.925 ;
        RECT 548.595 3.235 548.925 3.565 ;
        RECT 548.595 1.875 548.925 2.205 ;
        RECT 548.595 0.515 548.925 0.845 ;
        RECT 548.6 -8.32 548.92 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 549.955 15.475 550.285 15.805 ;
        RECT 549.955 10.035 550.285 10.365 ;
        RECT 549.955 8.675 550.285 9.005 ;
        RECT 549.955 7.315 550.285 7.645 ;
        RECT 549.955 5.955 550.285 6.285 ;
        RECT 549.955 4.595 550.285 4.925 ;
        RECT 549.955 3.235 550.285 3.565 ;
        RECT 549.955 1.875 550.285 2.205 ;
        RECT 549.955 0.515 550.285 0.845 ;
        RECT 549.96 -8.32 550.28 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 551.315 15.475 551.645 15.805 ;
        RECT 551.315 10.035 551.645 10.365 ;
        RECT 551.315 8.675 551.645 9.005 ;
        RECT 551.315 7.315 551.645 7.645 ;
        RECT 551.315 5.955 551.645 6.285 ;
        RECT 551.315 4.595 551.645 4.925 ;
        RECT 551.315 3.235 551.645 3.565 ;
        RECT 551.315 1.875 551.645 2.205 ;
        RECT 551.315 0.515 551.645 0.845 ;
        RECT 551.32 -8.32 551.64 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 552.675 15.475 553.005 15.805 ;
        RECT 552.675 10.035 553.005 10.365 ;
        RECT 552.675 8.675 553.005 9.005 ;
        RECT 552.675 7.315 553.005 7.645 ;
        RECT 552.675 5.955 553.005 6.285 ;
        RECT 552.675 4.595 553.005 4.925 ;
        RECT 552.675 3.235 553.005 3.565 ;
        RECT 552.675 1.875 553.005 2.205 ;
        RECT 552.675 0.515 553.005 0.845 ;
        RECT 552.68 -8.32 553 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 554.035 15.475 554.365 15.805 ;
        RECT 554.035 10.035 554.365 10.365 ;
        RECT 554.035 8.675 554.365 9.005 ;
        RECT 554.035 7.315 554.365 7.645 ;
        RECT 554.035 5.955 554.365 6.285 ;
        RECT 554.035 4.595 554.365 4.925 ;
        RECT 554.035 3.235 554.365 3.565 ;
        RECT 554.035 1.875 554.365 2.205 ;
        RECT 554.035 0.515 554.365 0.845 ;
        RECT 554.04 -8.32 554.36 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 555.395 15.475 555.725 15.805 ;
        RECT 555.395 11.395 555.725 11.725 ;
        RECT 555.395 10.035 555.725 10.365 ;
        RECT 555.395 8.675 555.725 9.005 ;
        RECT 555.395 7.315 555.725 7.645 ;
        RECT 555.395 5.955 555.725 6.285 ;
        RECT 555.395 4.595 555.725 4.925 ;
        RECT 555.395 3.235 555.725 3.565 ;
        RECT 555.395 1.875 555.725 2.205 ;
        RECT 555.395 0.515 555.725 0.845 ;
        RECT 555.4 -8.32 555.72 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 556.755 15.475 557.085 15.805 ;
        RECT 556.755 11.395 557.085 11.725 ;
        RECT 556.755 10.035 557.085 10.365 ;
        RECT 556.755 8.675 557.085 9.005 ;
        RECT 556.755 7.315 557.085 7.645 ;
        RECT 556.755 5.955 557.085 6.285 ;
        RECT 556.755 4.595 557.085 4.925 ;
        RECT 556.755 3.235 557.085 3.565 ;
        RECT 556.755 1.875 557.085 2.205 ;
        RECT 556.755 0.515 557.085 0.845 ;
        RECT 556.76 -8.32 557.08 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 558.115 15.475 558.445 15.805 ;
        RECT 558.115 11.395 558.445 11.725 ;
        RECT 558.115 10.035 558.445 10.365 ;
        RECT 558.115 8.675 558.445 9.005 ;
        RECT 558.115 7.315 558.445 7.645 ;
        RECT 558.115 5.955 558.445 6.285 ;
        RECT 558.115 4.595 558.445 4.925 ;
        RECT 558.115 3.235 558.445 3.565 ;
        RECT 558.115 1.875 558.445 2.205 ;
        RECT 558.115 0.515 558.445 0.845 ;
        RECT 558.12 -8.32 558.44 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 559.475 15.475 559.805 15.805 ;
        RECT 559.475 10.035 559.805 10.365 ;
        RECT 559.475 8.675 559.805 9.005 ;
        RECT 559.475 7.315 559.805 7.645 ;
        RECT 559.475 5.955 559.805 6.285 ;
        RECT 559.475 4.595 559.805 4.925 ;
        RECT 559.475 3.235 559.805 3.565 ;
        RECT 559.475 1.875 559.805 2.205 ;
        RECT 559.475 0.515 559.805 0.845 ;
        RECT 559.48 -8.32 559.8 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 560.835 15.475 561.165 15.805 ;
        RECT 560.835 10.035 561.165 10.365 ;
        RECT 560.835 8.675 561.165 9.005 ;
        RECT 560.835 7.315 561.165 7.645 ;
        RECT 560.835 5.955 561.165 6.285 ;
        RECT 560.835 4.595 561.165 4.925 ;
        RECT 560.835 3.235 561.165 3.565 ;
        RECT 560.835 1.875 561.165 2.205 ;
        RECT 560.835 0.515 561.165 0.845 ;
        RECT 560.84 -8.32 561.16 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 562.195 15.475 562.525 15.805 ;
        RECT 562.195 10.035 562.525 10.365 ;
        RECT 562.195 8.675 562.525 9.005 ;
        RECT 562.195 7.315 562.525 7.645 ;
        RECT 562.195 5.955 562.525 6.285 ;
        RECT 562.195 4.595 562.525 4.925 ;
        RECT 562.195 3.235 562.525 3.565 ;
        RECT 562.195 1.875 562.525 2.205 ;
        RECT 562.195 0.515 562.525 0.845 ;
        RECT 562.2 -8.32 562.52 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 563.555 15.475 563.885 15.805 ;
        RECT 563.555 10.035 563.885 10.365 ;
        RECT 563.555 8.675 563.885 9.005 ;
        RECT 563.555 7.315 563.885 7.645 ;
        RECT 563.555 5.955 563.885 6.285 ;
        RECT 563.555 4.595 563.885 4.925 ;
        RECT 563.555 3.235 563.885 3.565 ;
        RECT 563.555 1.875 563.885 2.205 ;
        RECT 563.555 0.515 563.885 0.845 ;
        RECT 563.56 -8.32 563.88 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 564.915 15.475 565.245 15.805 ;
        RECT 564.915 10.035 565.245 10.365 ;
        RECT 564.915 8.675 565.245 9.005 ;
        RECT 564.915 7.315 565.245 7.645 ;
        RECT 564.915 5.955 565.245 6.285 ;
        RECT 564.915 4.595 565.245 4.925 ;
        RECT 564.915 3.235 565.245 3.565 ;
        RECT 564.915 1.875 565.245 2.205 ;
        RECT 564.915 0.515 565.245 0.845 ;
        RECT 564.92 -8.32 565.24 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 566.275 15.475 566.605 15.805 ;
        RECT 566.275 10.035 566.605 10.365 ;
        RECT 566.275 8.675 566.605 9.005 ;
        RECT 566.275 7.315 566.605 7.645 ;
        RECT 566.275 5.955 566.605 6.285 ;
        RECT 566.275 4.595 566.605 4.925 ;
        RECT 566.275 3.235 566.605 3.565 ;
        RECT 566.275 1.875 566.605 2.205 ;
        RECT 566.275 0.515 566.605 0.845 ;
        RECT 566.28 -8.32 566.6 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 567.635 15.475 567.965 15.805 ;
        RECT 567.635 11.395 567.965 11.725 ;
        RECT 567.635 10.035 567.965 10.365 ;
        RECT 567.635 8.675 567.965 9.005 ;
        RECT 567.635 7.315 567.965 7.645 ;
        RECT 567.635 5.955 567.965 6.285 ;
        RECT 567.635 4.595 567.965 4.925 ;
        RECT 567.635 3.235 567.965 3.565 ;
        RECT 567.635 1.875 567.965 2.205 ;
        RECT 567.635 0.515 567.965 0.845 ;
        RECT 567.64 -8.32 567.96 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 568.995 15.475 569.325 15.805 ;
        RECT 568.995 11.395 569.325 11.725 ;
        RECT 568.995 10.035 569.325 10.365 ;
        RECT 568.995 8.675 569.325 9.005 ;
        RECT 568.995 7.315 569.325 7.645 ;
        RECT 568.995 5.955 569.325 6.285 ;
        RECT 568.995 4.595 569.325 4.925 ;
        RECT 568.995 3.235 569.325 3.565 ;
        RECT 568.995 1.875 569.325 2.205 ;
        RECT 568.995 0.515 569.325 0.845 ;
        RECT 569 -8.32 569.32 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 570.355 15.475 570.685 15.805 ;
        RECT 570.355 11.395 570.685 11.725 ;
        RECT 570.355 10.035 570.685 10.365 ;
        RECT 570.355 8.675 570.685 9.005 ;
        RECT 570.355 7.315 570.685 7.645 ;
        RECT 570.355 5.955 570.685 6.285 ;
        RECT 570.355 4.595 570.685 4.925 ;
        RECT 570.355 3.235 570.685 3.565 ;
        RECT 570.355 1.875 570.685 2.205 ;
        RECT 570.355 0.515 570.685 0.845 ;
        RECT 570.36 -8.32 570.68 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 571.715 15.475 572.045 15.805 ;
        RECT 571.715 10.035 572.045 10.365 ;
        RECT 571.715 8.675 572.045 9.005 ;
        RECT 571.715 7.315 572.045 7.645 ;
        RECT 571.715 5.955 572.045 6.285 ;
        RECT 571.715 4.595 572.045 4.925 ;
        RECT 571.715 3.235 572.045 3.565 ;
        RECT 571.715 1.875 572.045 2.205 ;
        RECT 571.715 0.515 572.045 0.845 ;
        RECT 571.72 -8.32 572.04 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 573.075 15.475 573.405 15.805 ;
        RECT 573.075 10.035 573.405 10.365 ;
        RECT 573.075 8.675 573.405 9.005 ;
        RECT 573.075 7.315 573.405 7.645 ;
        RECT 573.075 5.955 573.405 6.285 ;
        RECT 573.075 4.595 573.405 4.925 ;
        RECT 573.075 3.235 573.405 3.565 ;
        RECT 573.075 1.875 573.405 2.205 ;
        RECT 573.075 0.515 573.405 0.845 ;
        RECT 573.08 -8.32 573.4 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 574.435 15.475 574.765 15.805 ;
        RECT 574.435 10.035 574.765 10.365 ;
        RECT 574.435 8.675 574.765 9.005 ;
        RECT 574.435 7.315 574.765 7.645 ;
        RECT 574.435 5.955 574.765 6.285 ;
        RECT 574.435 4.595 574.765 4.925 ;
        RECT 574.435 3.235 574.765 3.565 ;
        RECT 574.435 1.875 574.765 2.205 ;
        RECT 574.435 0.515 574.765 0.845 ;
        RECT 574.44 -8.32 574.76 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 575.795 15.475 576.125 15.805 ;
        RECT 575.795 10.035 576.125 10.365 ;
        RECT 575.795 8.675 576.125 9.005 ;
        RECT 575.795 7.315 576.125 7.645 ;
        RECT 575.795 5.955 576.125 6.285 ;
        RECT 575.795 4.595 576.125 4.925 ;
        RECT 575.795 3.235 576.125 3.565 ;
        RECT 575.795 1.875 576.125 2.205 ;
        RECT 575.795 0.515 576.125 0.845 ;
        RECT 575.8 -8.32 576.12 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 577.155 15.475 577.485 15.805 ;
        RECT 577.155 10.035 577.485 10.365 ;
        RECT 577.155 8.675 577.485 9.005 ;
        RECT 577.155 7.315 577.485 7.645 ;
        RECT 577.155 5.955 577.485 6.285 ;
        RECT 577.155 4.595 577.485 4.925 ;
        RECT 577.155 3.235 577.485 3.565 ;
        RECT 577.155 1.875 577.485 2.205 ;
        RECT 577.155 0.515 577.485 0.845 ;
        RECT 577.16 -8.32 577.48 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 578.515 15.475 578.845 15.805 ;
        RECT 578.515 10.035 578.845 10.365 ;
        RECT 578.515 8.675 578.845 9.005 ;
        RECT 578.515 7.315 578.845 7.645 ;
        RECT 578.515 5.955 578.845 6.285 ;
        RECT 578.515 4.595 578.845 4.925 ;
        RECT 578.515 3.235 578.845 3.565 ;
        RECT 578.515 1.875 578.845 2.205 ;
        RECT 578.515 0.515 578.845 0.845 ;
        RECT 578.52 -8.32 578.84 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 579.875 15.475 580.205 15.805 ;
        RECT 579.875 11.395 580.205 11.725 ;
        RECT 579.875 10.035 580.205 10.365 ;
        RECT 579.875 8.675 580.205 9.005 ;
        RECT 579.875 7.315 580.205 7.645 ;
        RECT 579.875 5.955 580.205 6.285 ;
        RECT 579.875 4.595 580.205 4.925 ;
        RECT 579.875 3.235 580.205 3.565 ;
        RECT 579.875 1.875 580.205 2.205 ;
        RECT 579.875 0.515 580.205 0.845 ;
        RECT 579.88 -8.32 580.2 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 581.235 15.475 581.565 15.805 ;
        RECT 581.235 11.395 581.565 11.725 ;
        RECT 581.235 10.035 581.565 10.365 ;
        RECT 581.235 8.675 581.565 9.005 ;
        RECT 581.235 7.315 581.565 7.645 ;
        RECT 581.235 5.955 581.565 6.285 ;
        RECT 581.235 4.595 581.565 4.925 ;
        RECT 581.235 3.235 581.565 3.565 ;
        RECT 581.235 1.875 581.565 2.205 ;
        RECT 581.235 0.515 581.565 0.845 ;
        RECT 581.24 -8.32 581.56 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 582.595 15.475 582.925 15.805 ;
        RECT 582.595 11.395 582.925 11.725 ;
        RECT 582.595 10.035 582.925 10.365 ;
        RECT 582.595 8.675 582.925 9.005 ;
        RECT 582.595 7.315 582.925 7.645 ;
        RECT 582.595 5.955 582.925 6.285 ;
        RECT 582.595 4.595 582.925 4.925 ;
        RECT 582.595 3.235 582.925 3.565 ;
        RECT 582.595 1.875 582.925 2.205 ;
        RECT 582.595 0.515 582.925 0.845 ;
        RECT 582.6 -8.32 582.92 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 583.955 15.475 584.285 15.805 ;
        RECT 583.955 10.035 584.285 10.365 ;
        RECT 583.955 8.675 584.285 9.005 ;
        RECT 583.955 7.315 584.285 7.645 ;
        RECT 583.955 5.955 584.285 6.285 ;
        RECT 583.955 4.595 584.285 4.925 ;
        RECT 583.955 3.235 584.285 3.565 ;
        RECT 583.955 1.875 584.285 2.205 ;
        RECT 583.955 0.515 584.285 0.845 ;
        RECT 583.96 -8.32 584.28 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 585.315 15.475 585.645 15.805 ;
        RECT 585.315 10.035 585.645 10.365 ;
        RECT 585.315 8.675 585.645 9.005 ;
        RECT 585.315 7.315 585.645 7.645 ;
        RECT 585.315 5.955 585.645 6.285 ;
        RECT 585.315 4.595 585.645 4.925 ;
        RECT 585.315 3.235 585.645 3.565 ;
        RECT 585.315 1.875 585.645 2.205 ;
        RECT 585.315 0.515 585.645 0.845 ;
        RECT 585.32 -8.32 585.64 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 586.675 15.475 587.005 15.805 ;
        RECT 586.675 10.035 587.005 10.365 ;
        RECT 586.675 8.675 587.005 9.005 ;
        RECT 586.675 7.315 587.005 7.645 ;
        RECT 586.675 5.955 587.005 6.285 ;
        RECT 586.675 4.595 587.005 4.925 ;
        RECT 586.675 3.235 587.005 3.565 ;
        RECT 586.675 1.875 587.005 2.205 ;
        RECT 586.675 0.515 587.005 0.845 ;
        RECT 586.68 -8.32 587 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 588.035 15.475 588.365 15.805 ;
        RECT 588.035 10.035 588.365 10.365 ;
        RECT 588.035 8.675 588.365 9.005 ;
        RECT 588.035 7.315 588.365 7.645 ;
        RECT 588.035 5.955 588.365 6.285 ;
        RECT 588.035 4.595 588.365 4.925 ;
        RECT 588.035 3.235 588.365 3.565 ;
        RECT 588.035 1.875 588.365 2.205 ;
        RECT 588.035 0.515 588.365 0.845 ;
        RECT 588.04 -8.32 588.36 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 589.395 15.475 589.725 15.805 ;
        RECT 589.395 10.035 589.725 10.365 ;
        RECT 589.395 8.675 589.725 9.005 ;
        RECT 589.395 7.315 589.725 7.645 ;
        RECT 589.395 5.955 589.725 6.285 ;
        RECT 589.395 4.595 589.725 4.925 ;
        RECT 589.395 3.235 589.725 3.565 ;
        RECT 589.395 1.875 589.725 2.205 ;
        RECT 589.395 0.515 589.725 0.845 ;
        RECT 589.4 -8.32 589.72 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 590.755 15.475 591.085 15.805 ;
        RECT 590.755 10.035 591.085 10.365 ;
        RECT 590.755 8.675 591.085 9.005 ;
        RECT 590.755 7.315 591.085 7.645 ;
        RECT 590.755 5.955 591.085 6.285 ;
        RECT 590.755 4.595 591.085 4.925 ;
        RECT 590.755 3.235 591.085 3.565 ;
        RECT 590.755 1.875 591.085 2.205 ;
        RECT 590.755 0.515 591.085 0.845 ;
        RECT 590.76 -8.32 591.08 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 592.115 15.475 592.445 15.805 ;
        RECT 592.115 11.395 592.445 11.725 ;
        RECT 592.115 10.035 592.445 10.365 ;
        RECT 592.115 8.675 592.445 9.005 ;
        RECT 592.115 7.315 592.445 7.645 ;
        RECT 592.115 5.955 592.445 6.285 ;
        RECT 592.115 4.595 592.445 4.925 ;
        RECT 592.115 3.235 592.445 3.565 ;
        RECT 592.115 1.875 592.445 2.205 ;
        RECT 592.115 0.515 592.445 0.845 ;
        RECT 592.12 -8.32 592.44 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 593.475 15.475 593.805 15.805 ;
        RECT 593.475 11.395 593.805 11.725 ;
        RECT 593.475 10.035 593.805 10.365 ;
        RECT 593.475 8.675 593.805 9.005 ;
        RECT 593.475 7.315 593.805 7.645 ;
        RECT 593.475 5.955 593.805 6.285 ;
        RECT 593.475 4.595 593.805 4.925 ;
        RECT 593.475 3.235 593.805 3.565 ;
        RECT 593.475 1.875 593.805 2.205 ;
        RECT 593.475 0.515 593.805 0.845 ;
        RECT 593.48 -8.32 593.8 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 594.835 15.475 595.165 15.805 ;
        RECT 594.835 11.395 595.165 11.725 ;
        RECT 594.835 10.035 595.165 10.365 ;
        RECT 594.835 8.675 595.165 9.005 ;
        RECT 594.835 7.315 595.165 7.645 ;
        RECT 594.835 5.955 595.165 6.285 ;
        RECT 594.835 4.595 595.165 4.925 ;
        RECT 594.835 3.235 595.165 3.565 ;
        RECT 594.835 1.875 595.165 2.205 ;
        RECT 594.835 0.515 595.165 0.845 ;
        RECT 594.84 -8.32 595.16 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 596.195 15.475 596.525 15.805 ;
        RECT 596.195 10.035 596.525 10.365 ;
        RECT 596.195 8.675 596.525 9.005 ;
        RECT 596.195 7.315 596.525 7.645 ;
        RECT 596.195 5.955 596.525 6.285 ;
        RECT 596.195 4.595 596.525 4.925 ;
        RECT 596.195 3.235 596.525 3.565 ;
        RECT 596.195 1.875 596.525 2.205 ;
        RECT 596.195 0.515 596.525 0.845 ;
        RECT 596.2 -8.32 596.52 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 597.555 15.475 597.885 15.805 ;
        RECT 597.555 10.035 597.885 10.365 ;
        RECT 597.555 8.675 597.885 9.005 ;
        RECT 597.555 7.315 597.885 7.645 ;
        RECT 597.555 5.955 597.885 6.285 ;
        RECT 597.555 4.595 597.885 4.925 ;
        RECT 597.555 3.235 597.885 3.565 ;
        RECT 597.555 1.875 597.885 2.205 ;
        RECT 597.555 0.515 597.885 0.845 ;
        RECT 597.56 -8.32 597.88 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 598.915 15.475 599.245 15.805 ;
        RECT 598.915 10.035 599.245 10.365 ;
        RECT 598.915 8.675 599.245 9.005 ;
        RECT 598.915 7.315 599.245 7.645 ;
        RECT 598.915 5.955 599.245 6.285 ;
        RECT 598.915 4.595 599.245 4.925 ;
        RECT 598.915 3.235 599.245 3.565 ;
        RECT 598.915 1.875 599.245 2.205 ;
        RECT 598.915 0.515 599.245 0.845 ;
        RECT 598.92 -8.32 599.24 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 600.275 15.475 600.605 15.805 ;
        RECT 600.275 10.035 600.605 10.365 ;
        RECT 600.275 8.675 600.605 9.005 ;
        RECT 600.275 7.315 600.605 7.645 ;
        RECT 600.275 5.955 600.605 6.285 ;
        RECT 600.275 4.595 600.605 4.925 ;
        RECT 600.275 3.235 600.605 3.565 ;
        RECT 600.275 1.875 600.605 2.205 ;
        RECT 600.275 0.515 600.605 0.845 ;
        RECT 600.28 -8.32 600.6 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 601.635 15.475 601.965 15.805 ;
        RECT 601.635 10.035 601.965 10.365 ;
        RECT 601.635 8.675 601.965 9.005 ;
        RECT 601.635 7.315 601.965 7.645 ;
        RECT 601.635 5.955 601.965 6.285 ;
        RECT 601.635 4.595 601.965 4.925 ;
        RECT 601.635 3.235 601.965 3.565 ;
        RECT 601.635 1.875 601.965 2.205 ;
        RECT 601.635 0.515 601.965 0.845 ;
        RECT 601.64 -8.32 601.96 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 602.995 15.475 603.325 15.805 ;
        RECT 602.995 11.395 603.325 11.725 ;
        RECT 602.995 10.035 603.325 10.365 ;
        RECT 602.995 8.675 603.325 9.005 ;
        RECT 602.995 7.315 603.325 7.645 ;
        RECT 602.995 5.955 603.325 6.285 ;
        RECT 602.995 4.595 603.325 4.925 ;
        RECT 602.995 3.235 603.325 3.565 ;
        RECT 602.995 1.875 603.325 2.205 ;
        RECT 602.995 0.515 603.325 0.845 ;
        RECT 603 -8.32 603.32 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 604.355 15.475 604.685 15.805 ;
        RECT 604.355 11.395 604.685 11.725 ;
        RECT 604.355 10.035 604.685 10.365 ;
        RECT 604.355 8.675 604.685 9.005 ;
        RECT 604.355 7.315 604.685 7.645 ;
        RECT 604.355 5.955 604.685 6.285 ;
        RECT 604.355 4.595 604.685 4.925 ;
        RECT 604.355 3.235 604.685 3.565 ;
        RECT 604.355 1.875 604.685 2.205 ;
        RECT 604.355 0.515 604.685 0.845 ;
        RECT 604.36 -8.32 604.68 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 605.715 15.475 606.045 15.805 ;
        RECT 605.715 11.395 606.045 11.725 ;
        RECT 605.715 10.035 606.045 10.365 ;
        RECT 605.715 8.675 606.045 9.005 ;
        RECT 605.715 7.315 606.045 7.645 ;
        RECT 605.715 5.955 606.045 6.285 ;
        RECT 605.715 4.595 606.045 4.925 ;
        RECT 605.715 3.235 606.045 3.565 ;
        RECT 605.715 1.875 606.045 2.205 ;
        RECT 605.715 0.515 606.045 0.845 ;
        RECT 605.72 -8.32 606.04 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 607.075 15.475 607.405 15.805 ;
        RECT 607.075 10.035 607.405 10.365 ;
        RECT 607.075 8.675 607.405 9.005 ;
        RECT 607.075 7.315 607.405 7.645 ;
        RECT 607.075 5.955 607.405 6.285 ;
        RECT 607.075 4.595 607.405 4.925 ;
        RECT 607.075 3.235 607.405 3.565 ;
        RECT 607.075 1.875 607.405 2.205 ;
        RECT 607.075 0.515 607.405 0.845 ;
        RECT 607.08 -8.32 607.4 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 608.435 15.475 608.765 15.805 ;
        RECT 608.435 10.035 608.765 10.365 ;
        RECT 608.435 8.675 608.765 9.005 ;
        RECT 608.435 7.315 608.765 7.645 ;
        RECT 608.435 5.955 608.765 6.285 ;
        RECT 608.435 4.595 608.765 4.925 ;
        RECT 608.435 3.235 608.765 3.565 ;
        RECT 608.435 1.875 608.765 2.205 ;
        RECT 608.435 0.515 608.765 0.845 ;
        RECT 608.44 -8.32 608.76 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 609.795 15.475 610.125 15.805 ;
        RECT 609.795 10.035 610.125 10.365 ;
        RECT 609.795 8.675 610.125 9.005 ;
        RECT 609.795 7.315 610.125 7.645 ;
        RECT 609.795 5.955 610.125 6.285 ;
        RECT 609.795 4.595 610.125 4.925 ;
        RECT 609.795 3.235 610.125 3.565 ;
        RECT 609.795 1.875 610.125 2.205 ;
        RECT 609.795 0.515 610.125 0.845 ;
        RECT 609.8 -8.32 610.12 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 611.155 15.475 611.485 15.805 ;
        RECT 611.155 10.035 611.485 10.365 ;
        RECT 611.155 8.675 611.485 9.005 ;
        RECT 611.155 7.315 611.485 7.645 ;
        RECT 611.155 5.955 611.485 6.285 ;
        RECT 611.155 4.595 611.485 4.925 ;
        RECT 611.155 3.235 611.485 3.565 ;
        RECT 611.155 1.875 611.485 2.205 ;
        RECT 611.155 0.515 611.485 0.845 ;
        RECT 611.16 -8.32 611.48 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 612.515 15.475 612.845 15.805 ;
        RECT 612.515 10.035 612.845 10.365 ;
        RECT 612.515 8.675 612.845 9.005 ;
        RECT 612.515 7.315 612.845 7.645 ;
        RECT 612.515 5.955 612.845 6.285 ;
        RECT 612.515 4.595 612.845 4.925 ;
        RECT 612.515 3.235 612.845 3.565 ;
        RECT 612.515 1.875 612.845 2.205 ;
        RECT 612.515 0.515 612.845 0.845 ;
        RECT 612.52 -8.32 612.84 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 613.875 15.475 614.205 15.805 ;
        RECT 613.875 10.035 614.205 10.365 ;
        RECT 613.875 8.675 614.205 9.005 ;
        RECT 613.875 7.315 614.205 7.645 ;
        RECT 613.875 5.955 614.205 6.285 ;
        RECT 613.875 4.595 614.205 4.925 ;
        RECT 613.875 3.235 614.205 3.565 ;
        RECT 613.875 1.875 614.205 2.205 ;
        RECT 613.875 0.515 614.205 0.845 ;
        RECT 613.88 -8.32 614.2 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 615.235 15.475 615.565 15.805 ;
        RECT 615.235 11.395 615.565 11.725 ;
        RECT 615.235 10.035 615.565 10.365 ;
        RECT 615.235 8.675 615.565 9.005 ;
        RECT 615.235 7.315 615.565 7.645 ;
        RECT 615.235 5.955 615.565 6.285 ;
        RECT 615.235 4.595 615.565 4.925 ;
        RECT 615.235 3.235 615.565 3.565 ;
        RECT 615.235 1.875 615.565 2.205 ;
        RECT 615.235 0.515 615.565 0.845 ;
        RECT 615.24 -8.32 615.56 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 616.595 15.475 616.925 15.805 ;
        RECT 616.595 11.395 616.925 11.725 ;
        RECT 616.595 10.035 616.925 10.365 ;
        RECT 616.595 8.675 616.925 9.005 ;
        RECT 616.595 7.315 616.925 7.645 ;
        RECT 616.595 5.955 616.925 6.285 ;
        RECT 616.595 4.595 616.925 4.925 ;
        RECT 616.595 3.235 616.925 3.565 ;
        RECT 616.595 1.875 616.925 2.205 ;
        RECT 616.595 0.515 616.925 0.845 ;
        RECT 616.6 -8.32 616.92 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 617.955 15.475 618.285 15.805 ;
        RECT 617.955 11.395 618.285 11.725 ;
        RECT 617.955 10.035 618.285 10.365 ;
        RECT 617.955 8.675 618.285 9.005 ;
        RECT 617.955 7.315 618.285 7.645 ;
        RECT 617.955 5.955 618.285 6.285 ;
        RECT 617.955 4.595 618.285 4.925 ;
        RECT 617.955 3.235 618.285 3.565 ;
        RECT 617.955 1.875 618.285 2.205 ;
        RECT 617.955 0.515 618.285 0.845 ;
        RECT 617.96 -8.32 618.28 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 619.315 15.475 619.645 15.805 ;
        RECT 619.315 10.035 619.645 10.365 ;
        RECT 619.315 8.675 619.645 9.005 ;
        RECT 619.315 7.315 619.645 7.645 ;
        RECT 619.315 5.955 619.645 6.285 ;
        RECT 619.315 4.595 619.645 4.925 ;
        RECT 619.315 3.235 619.645 3.565 ;
        RECT 619.315 1.875 619.645 2.205 ;
        RECT 619.315 0.515 619.645 0.845 ;
        RECT 619.32 -8.32 619.64 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 620.675 15.475 621.005 15.805 ;
        RECT 620.675 10.035 621.005 10.365 ;
        RECT 620.675 8.675 621.005 9.005 ;
        RECT 620.675 7.315 621.005 7.645 ;
        RECT 620.675 5.955 621.005 6.285 ;
        RECT 620.675 4.595 621.005 4.925 ;
        RECT 620.675 3.235 621.005 3.565 ;
        RECT 620.675 1.875 621.005 2.205 ;
        RECT 620.675 0.515 621.005 0.845 ;
        RECT 620.68 -8.32 621 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 622.035 15.475 622.365 15.805 ;
        RECT 622.035 10.035 622.365 10.365 ;
        RECT 622.035 8.675 622.365 9.005 ;
        RECT 622.035 7.315 622.365 7.645 ;
        RECT 622.035 5.955 622.365 6.285 ;
        RECT 622.035 4.595 622.365 4.925 ;
        RECT 622.035 3.235 622.365 3.565 ;
        RECT 622.035 1.875 622.365 2.205 ;
        RECT 622.035 0.515 622.365 0.845 ;
        RECT 622.04 -8.32 622.36 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 623.395 15.475 623.725 15.805 ;
        RECT 623.395 10.035 623.725 10.365 ;
        RECT 623.395 8.675 623.725 9.005 ;
        RECT 623.395 7.315 623.725 7.645 ;
        RECT 623.395 5.955 623.725 6.285 ;
        RECT 623.395 4.595 623.725 4.925 ;
        RECT 623.395 3.235 623.725 3.565 ;
        RECT 623.395 1.875 623.725 2.205 ;
        RECT 623.395 0.515 623.725 0.845 ;
        RECT 623.4 -8.32 623.72 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 624.755 15.475 625.085 15.805 ;
        RECT 624.755 10.035 625.085 10.365 ;
        RECT 624.755 8.675 625.085 9.005 ;
        RECT 624.755 7.315 625.085 7.645 ;
        RECT 624.755 5.955 625.085 6.285 ;
        RECT 624.755 4.595 625.085 4.925 ;
        RECT 624.755 3.235 625.085 3.565 ;
        RECT 624.755 1.875 625.085 2.205 ;
        RECT 624.755 0.515 625.085 0.845 ;
        RECT 624.76 -8.32 625.08 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 626.115 15.475 626.445 15.805 ;
        RECT 626.115 10.035 626.445 10.365 ;
        RECT 626.115 8.675 626.445 9.005 ;
        RECT 626.115 7.315 626.445 7.645 ;
        RECT 626.115 5.955 626.445 6.285 ;
        RECT 626.115 4.595 626.445 4.925 ;
        RECT 626.115 3.235 626.445 3.565 ;
        RECT 626.115 1.875 626.445 2.205 ;
        RECT 626.115 0.515 626.445 0.845 ;
        RECT 626.12 -8.32 626.44 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 627.475 15.475 627.805 15.805 ;
        RECT 627.475 11.395 627.805 11.725 ;
        RECT 627.475 10.035 627.805 10.365 ;
        RECT 627.475 8.675 627.805 9.005 ;
        RECT 627.475 7.315 627.805 7.645 ;
        RECT 627.475 5.955 627.805 6.285 ;
        RECT 627.475 4.595 627.805 4.925 ;
        RECT 627.475 3.235 627.805 3.565 ;
        RECT 627.475 1.875 627.805 2.205 ;
        RECT 627.475 0.515 627.805 0.845 ;
        RECT 627.48 -8.32 627.8 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 628.835 15.475 629.165 15.805 ;
        RECT 628.835 11.395 629.165 11.725 ;
        RECT 628.835 10.035 629.165 10.365 ;
        RECT 628.835 8.675 629.165 9.005 ;
        RECT 628.835 7.315 629.165 7.645 ;
        RECT 628.835 5.955 629.165 6.285 ;
        RECT 628.835 4.595 629.165 4.925 ;
        RECT 628.835 3.235 629.165 3.565 ;
        RECT 628.835 1.875 629.165 2.205 ;
        RECT 628.835 0.515 629.165 0.845 ;
        RECT 628.84 -8.32 629.16 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 630.195 15.475 630.525 15.805 ;
        RECT 630.195 11.395 630.525 11.725 ;
        RECT 630.195 10.035 630.525 10.365 ;
        RECT 630.195 8.675 630.525 9.005 ;
        RECT 630.195 7.315 630.525 7.645 ;
        RECT 630.195 5.955 630.525 6.285 ;
        RECT 630.195 4.595 630.525 4.925 ;
        RECT 630.195 3.235 630.525 3.565 ;
        RECT 630.195 1.875 630.525 2.205 ;
        RECT 630.195 0.515 630.525 0.845 ;
        RECT 630.2 -8.32 630.52 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 631.555 15.475 631.885 15.805 ;
        RECT 631.555 10.035 631.885 10.365 ;
        RECT 631.555 8.675 631.885 9.005 ;
        RECT 631.555 7.315 631.885 7.645 ;
        RECT 631.555 5.955 631.885 6.285 ;
        RECT 631.555 4.595 631.885 4.925 ;
        RECT 631.555 3.235 631.885 3.565 ;
        RECT 631.555 1.875 631.885 2.205 ;
        RECT 631.555 0.515 631.885 0.845 ;
        RECT 631.56 -8.32 631.88 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 632.915 15.475 633.245 15.805 ;
        RECT 632.915 10.035 633.245 10.365 ;
        RECT 632.915 8.675 633.245 9.005 ;
        RECT 632.915 7.315 633.245 7.645 ;
        RECT 632.915 5.955 633.245 6.285 ;
        RECT 632.915 4.595 633.245 4.925 ;
        RECT 632.915 3.235 633.245 3.565 ;
        RECT 632.915 1.875 633.245 2.205 ;
        RECT 632.915 0.515 633.245 0.845 ;
        RECT 632.92 -8.32 633.24 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 634.275 15.475 634.605 15.805 ;
        RECT 634.275 10.035 634.605 10.365 ;
        RECT 634.275 8.675 634.605 9.005 ;
        RECT 634.275 7.315 634.605 7.645 ;
        RECT 634.275 5.955 634.605 6.285 ;
        RECT 634.275 4.595 634.605 4.925 ;
        RECT 634.275 3.235 634.605 3.565 ;
        RECT 634.275 1.875 634.605 2.205 ;
        RECT 634.275 0.515 634.605 0.845 ;
        RECT 634.28 -8.32 634.6 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 635.635 15.475 635.965 15.805 ;
        RECT 635.635 10.035 635.965 10.365 ;
        RECT 635.635 8.675 635.965 9.005 ;
        RECT 635.635 7.315 635.965 7.645 ;
        RECT 635.635 5.955 635.965 6.285 ;
        RECT 635.635 4.595 635.965 4.925 ;
        RECT 635.635 3.235 635.965 3.565 ;
        RECT 635.635 1.875 635.965 2.205 ;
        RECT 635.635 0.515 635.965 0.845 ;
        RECT 635.64 -8.32 635.96 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 636.995 15.475 637.325 15.805 ;
        RECT 636.995 10.035 637.325 10.365 ;
        RECT 636.995 8.675 637.325 9.005 ;
        RECT 636.995 7.315 637.325 7.645 ;
        RECT 636.995 5.955 637.325 6.285 ;
        RECT 636.995 4.595 637.325 4.925 ;
        RECT 636.995 3.235 637.325 3.565 ;
        RECT 636.995 1.875 637.325 2.205 ;
        RECT 636.995 0.515 637.325 0.845 ;
        RECT 637 -8.32 637.32 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 638.355 15.475 638.685 15.805 ;
        RECT 638.355 10.035 638.685 10.365 ;
        RECT 638.355 8.675 638.685 9.005 ;
        RECT 638.355 7.315 638.685 7.645 ;
        RECT 638.355 5.955 638.685 6.285 ;
        RECT 638.355 4.595 638.685 4.925 ;
        RECT 638.355 3.235 638.685 3.565 ;
        RECT 638.355 1.875 638.685 2.205 ;
        RECT 638.355 0.515 638.685 0.845 ;
        RECT 638.36 -8.32 638.68 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 639.715 3.235 640.045 3.565 ;
        RECT 639.715 1.875 640.045 2.205 ;
        RECT 639.715 0.515 640.045 0.845 ;
        RECT 639.72 -8.32 640.04 15.805 ;
        RECT 639.715 15.475 640.045 15.805 ;
        RECT 639.715 11.395 640.045 11.725 ;
        RECT 639.715 10.035 640.045 10.365 ;
        RECT 639.715 8.675 640.045 9.005 ;
        RECT 639.715 7.315 640.045 7.645 ;
        RECT 639.715 5.955 640.045 6.285 ;
        RECT 639.715 4.595 640.045 4.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 377.235 15.475 377.565 15.805 ;
        RECT 377.235 11.395 377.565 11.725 ;
        RECT 377.235 10.035 377.565 10.365 ;
        RECT 377.235 8.675 377.565 9.005 ;
        RECT 377.235 7.315 377.565 7.645 ;
        RECT 377.235 5.955 377.565 6.285 ;
        RECT 377.235 4.595 377.565 4.925 ;
        RECT 377.235 3.235 377.565 3.565 ;
        RECT 377.235 1.875 377.565 2.205 ;
        RECT 377.235 0.515 377.565 0.845 ;
        RECT 377.24 -8.32 377.56 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 378.595 15.475 378.925 15.805 ;
        RECT 378.595 11.395 378.925 11.725 ;
        RECT 378.595 10.035 378.925 10.365 ;
        RECT 378.595 8.675 378.925 9.005 ;
        RECT 378.595 7.315 378.925 7.645 ;
        RECT 378.595 5.955 378.925 6.285 ;
        RECT 378.595 4.595 378.925 4.925 ;
        RECT 378.595 3.235 378.925 3.565 ;
        RECT 378.595 1.875 378.925 2.205 ;
        RECT 378.595 0.515 378.925 0.845 ;
        RECT 378.6 -8.32 378.92 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 379.955 15.475 380.285 15.805 ;
        RECT 379.955 10.035 380.285 10.365 ;
        RECT 379.955 8.675 380.285 9.005 ;
        RECT 379.955 7.315 380.285 7.645 ;
        RECT 379.955 5.955 380.285 6.285 ;
        RECT 379.955 4.595 380.285 4.925 ;
        RECT 379.955 3.235 380.285 3.565 ;
        RECT 379.955 1.875 380.285 2.205 ;
        RECT 379.955 0.515 380.285 0.845 ;
        RECT 379.96 -8.32 380.28 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 381.315 15.475 381.645 15.805 ;
        RECT 381.315 10.035 381.645 10.365 ;
        RECT 381.315 8.675 381.645 9.005 ;
        RECT 381.315 7.315 381.645 7.645 ;
        RECT 381.315 5.955 381.645 6.285 ;
        RECT 381.315 4.595 381.645 4.925 ;
        RECT 381.315 3.235 381.645 3.565 ;
        RECT 381.315 1.875 381.645 2.205 ;
        RECT 381.315 0.515 381.645 0.845 ;
        RECT 381.32 -8.32 381.64 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 382.675 15.475 383.005 15.805 ;
        RECT 382.675 10.035 383.005 10.365 ;
        RECT 382.675 8.675 383.005 9.005 ;
        RECT 382.675 7.315 383.005 7.645 ;
        RECT 382.675 5.955 383.005 6.285 ;
        RECT 382.675 4.595 383.005 4.925 ;
        RECT 382.675 3.235 383.005 3.565 ;
        RECT 382.675 1.875 383.005 2.205 ;
        RECT 382.675 0.515 383.005 0.845 ;
        RECT 382.68 -8.32 383 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 384.035 15.475 384.365 15.805 ;
        RECT 384.035 10.035 384.365 10.365 ;
        RECT 384.035 8.675 384.365 9.005 ;
        RECT 384.035 7.315 384.365 7.645 ;
        RECT 384.035 5.955 384.365 6.285 ;
        RECT 384.035 4.595 384.365 4.925 ;
        RECT 384.035 3.235 384.365 3.565 ;
        RECT 384.035 1.875 384.365 2.205 ;
        RECT 384.035 0.515 384.365 0.845 ;
        RECT 384.04 -8.32 384.36 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 385.395 15.475 385.725 15.805 ;
        RECT 385.395 10.035 385.725 10.365 ;
        RECT 385.395 8.675 385.725 9.005 ;
        RECT 385.395 7.315 385.725 7.645 ;
        RECT 385.395 5.955 385.725 6.285 ;
        RECT 385.395 4.595 385.725 4.925 ;
        RECT 385.395 3.235 385.725 3.565 ;
        RECT 385.395 1.875 385.725 2.205 ;
        RECT 385.395 0.515 385.725 0.845 ;
        RECT 385.4 -8.32 385.72 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 386.755 15.475 387.085 15.805 ;
        RECT 386.755 10.035 387.085 10.365 ;
        RECT 386.755 8.675 387.085 9.005 ;
        RECT 386.755 7.315 387.085 7.645 ;
        RECT 386.755 5.955 387.085 6.285 ;
        RECT 386.755 4.595 387.085 4.925 ;
        RECT 386.755 3.235 387.085 3.565 ;
        RECT 386.755 1.875 387.085 2.205 ;
        RECT 386.755 0.515 387.085 0.845 ;
        RECT 386.76 -8.32 387.08 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 388.115 15.475 388.445 15.805 ;
        RECT 388.115 11.395 388.445 11.725 ;
        RECT 388.115 10.035 388.445 10.365 ;
        RECT 388.115 8.675 388.445 9.005 ;
        RECT 388.115 7.315 388.445 7.645 ;
        RECT 388.115 5.955 388.445 6.285 ;
        RECT 388.115 4.595 388.445 4.925 ;
        RECT 388.115 3.235 388.445 3.565 ;
        RECT 388.115 1.875 388.445 2.205 ;
        RECT 388.115 0.515 388.445 0.845 ;
        RECT 388.12 -8.32 388.44 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 389.475 15.475 389.805 15.805 ;
        RECT 389.475 11.395 389.805 11.725 ;
        RECT 389.475 10.035 389.805 10.365 ;
        RECT 389.475 8.675 389.805 9.005 ;
        RECT 389.475 7.315 389.805 7.645 ;
        RECT 389.475 5.955 389.805 6.285 ;
        RECT 389.475 4.595 389.805 4.925 ;
        RECT 389.475 3.235 389.805 3.565 ;
        RECT 389.475 1.875 389.805 2.205 ;
        RECT 389.475 0.515 389.805 0.845 ;
        RECT 389.48 -8.32 389.8 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 390.835 15.475 391.165 15.805 ;
        RECT 390.835 11.395 391.165 11.725 ;
        RECT 390.835 10.035 391.165 10.365 ;
        RECT 390.835 8.675 391.165 9.005 ;
        RECT 390.835 7.315 391.165 7.645 ;
        RECT 390.835 5.955 391.165 6.285 ;
        RECT 390.835 4.595 391.165 4.925 ;
        RECT 390.835 3.235 391.165 3.565 ;
        RECT 390.835 1.875 391.165 2.205 ;
        RECT 390.835 0.515 391.165 0.845 ;
        RECT 390.84 -8.32 391.16 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 392.195 15.475 392.525 15.805 ;
        RECT 392.195 10.035 392.525 10.365 ;
        RECT 392.195 8.675 392.525 9.005 ;
        RECT 392.195 7.315 392.525 7.645 ;
        RECT 392.195 5.955 392.525 6.285 ;
        RECT 392.195 4.595 392.525 4.925 ;
        RECT 392.195 3.235 392.525 3.565 ;
        RECT 392.195 1.875 392.525 2.205 ;
        RECT 392.195 0.515 392.525 0.845 ;
        RECT 392.2 -8.32 392.52 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 393.555 15.475 393.885 15.805 ;
        RECT 393.555 10.035 393.885 10.365 ;
        RECT 393.555 8.675 393.885 9.005 ;
        RECT 393.555 7.315 393.885 7.645 ;
        RECT 393.555 5.955 393.885 6.285 ;
        RECT 393.555 4.595 393.885 4.925 ;
        RECT 393.555 3.235 393.885 3.565 ;
        RECT 393.555 1.875 393.885 2.205 ;
        RECT 393.555 0.515 393.885 0.845 ;
        RECT 393.56 -8.32 393.88 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 394.915 15.475 395.245 15.805 ;
        RECT 394.915 10.035 395.245 10.365 ;
        RECT 394.915 8.675 395.245 9.005 ;
        RECT 394.915 7.315 395.245 7.645 ;
        RECT 394.915 5.955 395.245 6.285 ;
        RECT 394.915 4.595 395.245 4.925 ;
        RECT 394.915 3.235 395.245 3.565 ;
        RECT 394.915 1.875 395.245 2.205 ;
        RECT 394.915 0.515 395.245 0.845 ;
        RECT 394.92 -8.32 395.24 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 396.275 15.475 396.605 15.805 ;
        RECT 396.275 10.035 396.605 10.365 ;
        RECT 396.275 8.675 396.605 9.005 ;
        RECT 396.275 7.315 396.605 7.645 ;
        RECT 396.275 5.955 396.605 6.285 ;
        RECT 396.275 4.595 396.605 4.925 ;
        RECT 396.275 3.235 396.605 3.565 ;
        RECT 396.275 1.875 396.605 2.205 ;
        RECT 396.275 0.515 396.605 0.845 ;
        RECT 396.28 -8.32 396.6 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 397.635 15.475 397.965 15.805 ;
        RECT 397.635 10.035 397.965 10.365 ;
        RECT 397.635 8.675 397.965 9.005 ;
        RECT 397.635 7.315 397.965 7.645 ;
        RECT 397.635 5.955 397.965 6.285 ;
        RECT 397.635 4.595 397.965 4.925 ;
        RECT 397.635 3.235 397.965 3.565 ;
        RECT 397.635 1.875 397.965 2.205 ;
        RECT 397.635 0.515 397.965 0.845 ;
        RECT 397.64 -8.32 397.96 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 398.995 15.475 399.325 15.805 ;
        RECT 398.995 11.395 399.325 11.725 ;
        RECT 398.995 10.035 399.325 10.365 ;
        RECT 398.995 8.675 399.325 9.005 ;
        RECT 398.995 7.315 399.325 7.645 ;
        RECT 398.995 5.955 399.325 6.285 ;
        RECT 398.995 4.595 399.325 4.925 ;
        RECT 398.995 3.235 399.325 3.565 ;
        RECT 398.995 1.875 399.325 2.205 ;
        RECT 398.995 0.515 399.325 0.845 ;
        RECT 399 -8.32 399.32 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 400.355 15.475 400.685 15.805 ;
        RECT 400.355 11.395 400.685 11.725 ;
        RECT 400.355 10.035 400.685 10.365 ;
        RECT 400.355 8.675 400.685 9.005 ;
        RECT 400.355 7.315 400.685 7.645 ;
        RECT 400.355 5.955 400.685 6.285 ;
        RECT 400.355 4.595 400.685 4.925 ;
        RECT 400.355 3.235 400.685 3.565 ;
        RECT 400.355 1.875 400.685 2.205 ;
        RECT 400.355 0.515 400.685 0.845 ;
        RECT 400.36 -8.32 400.68 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 401.715 15.475 402.045 15.805 ;
        RECT 401.715 11.395 402.045 11.725 ;
        RECT 401.715 10.035 402.045 10.365 ;
        RECT 401.715 8.675 402.045 9.005 ;
        RECT 401.715 7.315 402.045 7.645 ;
        RECT 401.715 5.955 402.045 6.285 ;
        RECT 401.715 4.595 402.045 4.925 ;
        RECT 401.715 3.235 402.045 3.565 ;
        RECT 401.715 1.875 402.045 2.205 ;
        RECT 401.715 0.515 402.045 0.845 ;
        RECT 401.72 -8.32 402.04 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 403.075 15.475 403.405 15.805 ;
        RECT 403.075 10.035 403.405 10.365 ;
        RECT 403.075 8.675 403.405 9.005 ;
        RECT 403.075 7.315 403.405 7.645 ;
        RECT 403.075 5.955 403.405 6.285 ;
        RECT 403.075 4.595 403.405 4.925 ;
        RECT 403.075 3.235 403.405 3.565 ;
        RECT 403.075 1.875 403.405 2.205 ;
        RECT 403.075 0.515 403.405 0.845 ;
        RECT 403.08 -8.32 403.4 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 404.435 15.475 404.765 15.805 ;
        RECT 404.435 10.035 404.765 10.365 ;
        RECT 404.435 8.675 404.765 9.005 ;
        RECT 404.435 7.315 404.765 7.645 ;
        RECT 404.435 5.955 404.765 6.285 ;
        RECT 404.435 4.595 404.765 4.925 ;
        RECT 404.435 3.235 404.765 3.565 ;
        RECT 404.435 1.875 404.765 2.205 ;
        RECT 404.435 0.515 404.765 0.845 ;
        RECT 404.44 -8.32 404.76 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 405.795 15.475 406.125 15.805 ;
        RECT 405.795 10.035 406.125 10.365 ;
        RECT 405.795 8.675 406.125 9.005 ;
        RECT 405.795 7.315 406.125 7.645 ;
        RECT 405.795 5.955 406.125 6.285 ;
        RECT 405.795 4.595 406.125 4.925 ;
        RECT 405.795 3.235 406.125 3.565 ;
        RECT 405.795 1.875 406.125 2.205 ;
        RECT 405.795 0.515 406.125 0.845 ;
        RECT 405.8 -8.32 406.12 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 407.155 15.475 407.485 15.805 ;
        RECT 407.155 10.035 407.485 10.365 ;
        RECT 407.155 8.675 407.485 9.005 ;
        RECT 407.155 7.315 407.485 7.645 ;
        RECT 407.155 5.955 407.485 6.285 ;
        RECT 407.155 4.595 407.485 4.925 ;
        RECT 407.155 3.235 407.485 3.565 ;
        RECT 407.155 1.875 407.485 2.205 ;
        RECT 407.155 0.515 407.485 0.845 ;
        RECT 407.16 -8.32 407.48 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 408.515 15.475 408.845 15.805 ;
        RECT 408.515 10.035 408.845 10.365 ;
        RECT 408.515 8.675 408.845 9.005 ;
        RECT 408.515 7.315 408.845 7.645 ;
        RECT 408.515 5.955 408.845 6.285 ;
        RECT 408.515 4.595 408.845 4.925 ;
        RECT 408.515 3.235 408.845 3.565 ;
        RECT 408.515 1.875 408.845 2.205 ;
        RECT 408.515 0.515 408.845 0.845 ;
        RECT 408.52 -8.32 408.84 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 409.875 15.475 410.205 15.805 ;
        RECT 409.875 10.035 410.205 10.365 ;
        RECT 409.875 8.675 410.205 9.005 ;
        RECT 409.875 7.315 410.205 7.645 ;
        RECT 409.875 5.955 410.205 6.285 ;
        RECT 409.875 4.595 410.205 4.925 ;
        RECT 409.875 3.235 410.205 3.565 ;
        RECT 409.875 1.875 410.205 2.205 ;
        RECT 409.875 0.515 410.205 0.845 ;
        RECT 409.88 -8.32 410.2 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 411.235 15.475 411.565 15.805 ;
        RECT 411.235 11.395 411.565 11.725 ;
        RECT 411.235 10.035 411.565 10.365 ;
        RECT 411.235 8.675 411.565 9.005 ;
        RECT 411.235 7.315 411.565 7.645 ;
        RECT 411.235 5.955 411.565 6.285 ;
        RECT 411.235 4.595 411.565 4.925 ;
        RECT 411.235 3.235 411.565 3.565 ;
        RECT 411.235 1.875 411.565 2.205 ;
        RECT 411.235 0.515 411.565 0.845 ;
        RECT 411.24 -8.32 411.56 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 412.595 15.475 412.925 15.805 ;
        RECT 412.595 11.395 412.925 11.725 ;
        RECT 412.595 10.035 412.925 10.365 ;
        RECT 412.595 8.675 412.925 9.005 ;
        RECT 412.595 7.315 412.925 7.645 ;
        RECT 412.595 5.955 412.925 6.285 ;
        RECT 412.595 4.595 412.925 4.925 ;
        RECT 412.595 3.235 412.925 3.565 ;
        RECT 412.595 1.875 412.925 2.205 ;
        RECT 412.595 0.515 412.925 0.845 ;
        RECT 412.6 -8.32 412.92 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 413.955 15.475 414.285 15.805 ;
        RECT 413.955 11.395 414.285 11.725 ;
        RECT 413.955 10.035 414.285 10.365 ;
        RECT 413.955 8.675 414.285 9.005 ;
        RECT 413.955 7.315 414.285 7.645 ;
        RECT 413.955 5.955 414.285 6.285 ;
        RECT 413.955 4.595 414.285 4.925 ;
        RECT 413.955 3.235 414.285 3.565 ;
        RECT 413.955 1.875 414.285 2.205 ;
        RECT 413.955 0.515 414.285 0.845 ;
        RECT 413.96 -8.32 414.28 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 415.315 15.475 415.645 15.805 ;
        RECT 415.315 10.035 415.645 10.365 ;
        RECT 415.315 8.675 415.645 9.005 ;
        RECT 415.315 7.315 415.645 7.645 ;
        RECT 415.315 5.955 415.645 6.285 ;
        RECT 415.315 4.595 415.645 4.925 ;
        RECT 415.315 3.235 415.645 3.565 ;
        RECT 415.315 1.875 415.645 2.205 ;
        RECT 415.315 0.515 415.645 0.845 ;
        RECT 415.32 -8.32 415.64 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 416.675 15.475 417.005 15.805 ;
        RECT 416.675 10.035 417.005 10.365 ;
        RECT 416.675 8.675 417.005 9.005 ;
        RECT 416.675 7.315 417.005 7.645 ;
        RECT 416.675 5.955 417.005 6.285 ;
        RECT 416.675 4.595 417.005 4.925 ;
        RECT 416.675 3.235 417.005 3.565 ;
        RECT 416.675 1.875 417.005 2.205 ;
        RECT 416.675 0.515 417.005 0.845 ;
        RECT 416.68 -8.32 417 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 418.035 15.475 418.365 15.805 ;
        RECT 418.035 10.035 418.365 10.365 ;
        RECT 418.035 8.675 418.365 9.005 ;
        RECT 418.035 7.315 418.365 7.645 ;
        RECT 418.035 5.955 418.365 6.285 ;
        RECT 418.035 4.595 418.365 4.925 ;
        RECT 418.035 3.235 418.365 3.565 ;
        RECT 418.035 1.875 418.365 2.205 ;
        RECT 418.035 0.515 418.365 0.845 ;
        RECT 418.04 -8.32 418.36 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 419.395 15.475 419.725 15.805 ;
        RECT 419.395 10.035 419.725 10.365 ;
        RECT 419.395 8.675 419.725 9.005 ;
        RECT 419.395 7.315 419.725 7.645 ;
        RECT 419.395 5.955 419.725 6.285 ;
        RECT 419.395 4.595 419.725 4.925 ;
        RECT 419.395 3.235 419.725 3.565 ;
        RECT 419.395 1.875 419.725 2.205 ;
        RECT 419.395 0.515 419.725 0.845 ;
        RECT 419.4 -8.32 419.72 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 420.755 15.475 421.085 15.805 ;
        RECT 420.755 10.035 421.085 10.365 ;
        RECT 420.755 8.675 421.085 9.005 ;
        RECT 420.755 7.315 421.085 7.645 ;
        RECT 420.755 5.955 421.085 6.285 ;
        RECT 420.755 4.595 421.085 4.925 ;
        RECT 420.755 3.235 421.085 3.565 ;
        RECT 420.755 1.875 421.085 2.205 ;
        RECT 420.755 0.515 421.085 0.845 ;
        RECT 420.76 -8.32 421.08 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 422.115 15.475 422.445 15.805 ;
        RECT 422.115 10.035 422.445 10.365 ;
        RECT 422.115 8.675 422.445 9.005 ;
        RECT 422.115 7.315 422.445 7.645 ;
        RECT 422.115 5.955 422.445 6.285 ;
        RECT 422.115 4.595 422.445 4.925 ;
        RECT 422.115 3.235 422.445 3.565 ;
        RECT 422.115 1.875 422.445 2.205 ;
        RECT 422.115 0.515 422.445 0.845 ;
        RECT 422.12 -8.32 422.44 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 423.475 15.475 423.805 15.805 ;
        RECT 423.475 11.395 423.805 11.725 ;
        RECT 423.475 10.035 423.805 10.365 ;
        RECT 423.475 8.675 423.805 9.005 ;
        RECT 423.475 7.315 423.805 7.645 ;
        RECT 423.475 5.955 423.805 6.285 ;
        RECT 423.475 4.595 423.805 4.925 ;
        RECT 423.475 3.235 423.805 3.565 ;
        RECT 423.475 1.875 423.805 2.205 ;
        RECT 423.475 0.515 423.805 0.845 ;
        RECT 423.48 -8.32 423.8 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 424.835 15.475 425.165 15.805 ;
        RECT 424.835 11.395 425.165 11.725 ;
        RECT 424.835 10.035 425.165 10.365 ;
        RECT 424.835 8.675 425.165 9.005 ;
        RECT 424.835 7.315 425.165 7.645 ;
        RECT 424.835 5.955 425.165 6.285 ;
        RECT 424.835 4.595 425.165 4.925 ;
        RECT 424.835 3.235 425.165 3.565 ;
        RECT 424.835 1.875 425.165 2.205 ;
        RECT 424.835 0.515 425.165 0.845 ;
        RECT 424.84 -8.32 425.16 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 426.195 15.475 426.525 15.805 ;
        RECT 426.195 11.395 426.525 11.725 ;
        RECT 426.195 10.035 426.525 10.365 ;
        RECT 426.195 8.675 426.525 9.005 ;
        RECT 426.195 7.315 426.525 7.645 ;
        RECT 426.195 5.955 426.525 6.285 ;
        RECT 426.195 4.595 426.525 4.925 ;
        RECT 426.195 3.235 426.525 3.565 ;
        RECT 426.195 1.875 426.525 2.205 ;
        RECT 426.195 0.515 426.525 0.845 ;
        RECT 426.2 -8.32 426.52 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 427.555 15.475 427.885 15.805 ;
        RECT 427.555 10.035 427.885 10.365 ;
        RECT 427.555 8.675 427.885 9.005 ;
        RECT 427.555 7.315 427.885 7.645 ;
        RECT 427.555 5.955 427.885 6.285 ;
        RECT 427.555 4.595 427.885 4.925 ;
        RECT 427.555 3.235 427.885 3.565 ;
        RECT 427.555 1.875 427.885 2.205 ;
        RECT 427.555 0.515 427.885 0.845 ;
        RECT 427.56 -8.32 427.88 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 428.915 15.475 429.245 15.805 ;
        RECT 428.915 10.035 429.245 10.365 ;
        RECT 428.915 8.675 429.245 9.005 ;
        RECT 428.915 7.315 429.245 7.645 ;
        RECT 428.915 5.955 429.245 6.285 ;
        RECT 428.915 4.595 429.245 4.925 ;
        RECT 428.915 3.235 429.245 3.565 ;
        RECT 428.915 1.875 429.245 2.205 ;
        RECT 428.915 0.515 429.245 0.845 ;
        RECT 428.92 -8.32 429.24 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 430.275 15.475 430.605 15.805 ;
        RECT 430.275 10.035 430.605 10.365 ;
        RECT 430.275 8.675 430.605 9.005 ;
        RECT 430.275 7.315 430.605 7.645 ;
        RECT 430.275 5.955 430.605 6.285 ;
        RECT 430.275 4.595 430.605 4.925 ;
        RECT 430.275 3.235 430.605 3.565 ;
        RECT 430.275 1.875 430.605 2.205 ;
        RECT 430.275 0.515 430.605 0.845 ;
        RECT 430.28 -8.32 430.6 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 431.635 15.475 431.965 15.805 ;
        RECT 431.635 10.035 431.965 10.365 ;
        RECT 431.635 8.675 431.965 9.005 ;
        RECT 431.635 7.315 431.965 7.645 ;
        RECT 431.635 5.955 431.965 6.285 ;
        RECT 431.635 4.595 431.965 4.925 ;
        RECT 431.635 3.235 431.965 3.565 ;
        RECT 431.635 1.875 431.965 2.205 ;
        RECT 431.635 0.515 431.965 0.845 ;
        RECT 431.64 -8.32 431.96 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 432.995 15.475 433.325 15.805 ;
        RECT 432.995 10.035 433.325 10.365 ;
        RECT 432.995 8.675 433.325 9.005 ;
        RECT 432.995 7.315 433.325 7.645 ;
        RECT 432.995 5.955 433.325 6.285 ;
        RECT 432.995 4.595 433.325 4.925 ;
        RECT 432.995 3.235 433.325 3.565 ;
        RECT 432.995 1.875 433.325 2.205 ;
        RECT 432.995 0.515 433.325 0.845 ;
        RECT 433 -8.32 433.32 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 434.355 15.475 434.685 15.805 ;
        RECT 434.355 10.035 434.685 10.365 ;
        RECT 434.355 8.675 434.685 9.005 ;
        RECT 434.355 7.315 434.685 7.645 ;
        RECT 434.355 5.955 434.685 6.285 ;
        RECT 434.355 4.595 434.685 4.925 ;
        RECT 434.355 3.235 434.685 3.565 ;
        RECT 434.355 1.875 434.685 2.205 ;
        RECT 434.355 0.515 434.685 0.845 ;
        RECT 434.36 -8.32 434.68 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 435.715 15.475 436.045 15.805 ;
        RECT 435.715 11.395 436.045 11.725 ;
        RECT 435.715 10.035 436.045 10.365 ;
        RECT 435.715 8.675 436.045 9.005 ;
        RECT 435.715 7.315 436.045 7.645 ;
        RECT 435.715 5.955 436.045 6.285 ;
        RECT 435.715 4.595 436.045 4.925 ;
        RECT 435.715 3.235 436.045 3.565 ;
        RECT 435.715 1.875 436.045 2.205 ;
        RECT 435.715 0.515 436.045 0.845 ;
        RECT 435.72 -8.32 436.04 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 437.075 15.475 437.405 15.805 ;
        RECT 437.075 11.395 437.405 11.725 ;
        RECT 437.075 10.035 437.405 10.365 ;
        RECT 437.075 8.675 437.405 9.005 ;
        RECT 437.075 7.315 437.405 7.645 ;
        RECT 437.075 5.955 437.405 6.285 ;
        RECT 437.075 4.595 437.405 4.925 ;
        RECT 437.075 3.235 437.405 3.565 ;
        RECT 437.075 1.875 437.405 2.205 ;
        RECT 437.075 0.515 437.405 0.845 ;
        RECT 437.08 -8.32 437.4 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 438.435 15.475 438.765 15.805 ;
        RECT 438.435 11.395 438.765 11.725 ;
        RECT 438.435 10.035 438.765 10.365 ;
        RECT 438.435 8.675 438.765 9.005 ;
        RECT 438.435 7.315 438.765 7.645 ;
        RECT 438.435 5.955 438.765 6.285 ;
        RECT 438.435 4.595 438.765 4.925 ;
        RECT 438.435 3.235 438.765 3.565 ;
        RECT 438.435 1.875 438.765 2.205 ;
        RECT 438.435 0.515 438.765 0.845 ;
        RECT 438.44 -8.32 438.76 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 439.795 15.475 440.125 15.805 ;
        RECT 439.795 10.035 440.125 10.365 ;
        RECT 439.795 8.675 440.125 9.005 ;
        RECT 439.795 7.315 440.125 7.645 ;
        RECT 439.795 5.955 440.125 6.285 ;
        RECT 439.795 4.595 440.125 4.925 ;
        RECT 439.795 3.235 440.125 3.565 ;
        RECT 439.795 1.875 440.125 2.205 ;
        RECT 439.795 0.515 440.125 0.845 ;
        RECT 439.8 -8.32 440.12 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 441.155 15.475 441.485 15.805 ;
        RECT 441.155 10.035 441.485 10.365 ;
        RECT 441.155 8.675 441.485 9.005 ;
        RECT 441.155 7.315 441.485 7.645 ;
        RECT 441.155 5.955 441.485 6.285 ;
        RECT 441.155 4.595 441.485 4.925 ;
        RECT 441.155 3.235 441.485 3.565 ;
        RECT 441.155 1.875 441.485 2.205 ;
        RECT 441.155 0.515 441.485 0.845 ;
        RECT 441.16 -8.32 441.48 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 442.515 15.475 442.845 15.805 ;
        RECT 442.515 10.035 442.845 10.365 ;
        RECT 442.515 8.675 442.845 9.005 ;
        RECT 442.515 7.315 442.845 7.645 ;
        RECT 442.515 5.955 442.845 6.285 ;
        RECT 442.515 4.595 442.845 4.925 ;
        RECT 442.515 3.235 442.845 3.565 ;
        RECT 442.515 1.875 442.845 2.205 ;
        RECT 442.515 0.515 442.845 0.845 ;
        RECT 442.52 -8.32 442.84 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 443.875 15.475 444.205 15.805 ;
        RECT 443.875 10.035 444.205 10.365 ;
        RECT 443.875 8.675 444.205 9.005 ;
        RECT 443.875 7.315 444.205 7.645 ;
        RECT 443.875 5.955 444.205 6.285 ;
        RECT 443.875 4.595 444.205 4.925 ;
        RECT 443.875 3.235 444.205 3.565 ;
        RECT 443.875 1.875 444.205 2.205 ;
        RECT 443.875 0.515 444.205 0.845 ;
        RECT 443.88 -8.32 444.2 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 445.235 15.475 445.565 15.805 ;
        RECT 445.235 10.035 445.565 10.365 ;
        RECT 445.235 8.675 445.565 9.005 ;
        RECT 445.235 7.315 445.565 7.645 ;
        RECT 445.235 5.955 445.565 6.285 ;
        RECT 445.235 4.595 445.565 4.925 ;
        RECT 445.235 3.235 445.565 3.565 ;
        RECT 445.235 1.875 445.565 2.205 ;
        RECT 445.235 0.515 445.565 0.845 ;
        RECT 445.24 -8.32 445.56 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 446.595 15.475 446.925 15.805 ;
        RECT 446.595 10.035 446.925 10.365 ;
        RECT 446.595 8.675 446.925 9.005 ;
        RECT 446.595 7.315 446.925 7.645 ;
        RECT 446.595 5.955 446.925 6.285 ;
        RECT 446.595 4.595 446.925 4.925 ;
        RECT 446.595 3.235 446.925 3.565 ;
        RECT 446.595 1.875 446.925 2.205 ;
        RECT 446.595 0.515 446.925 0.845 ;
        RECT 446.6 -8.32 446.92 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 447.955 15.475 448.285 15.805 ;
        RECT 447.955 11.395 448.285 11.725 ;
        RECT 447.955 10.035 448.285 10.365 ;
        RECT 447.955 8.675 448.285 9.005 ;
        RECT 447.955 7.315 448.285 7.645 ;
        RECT 447.955 5.955 448.285 6.285 ;
        RECT 447.955 4.595 448.285 4.925 ;
        RECT 447.955 3.235 448.285 3.565 ;
        RECT 447.955 1.875 448.285 2.205 ;
        RECT 447.955 0.515 448.285 0.845 ;
        RECT 447.96 -8.32 448.28 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 449.315 15.475 449.645 15.805 ;
        RECT 449.315 11.395 449.645 11.725 ;
        RECT 449.315 10.035 449.645 10.365 ;
        RECT 449.315 8.675 449.645 9.005 ;
        RECT 449.315 7.315 449.645 7.645 ;
        RECT 449.315 5.955 449.645 6.285 ;
        RECT 449.315 4.595 449.645 4.925 ;
        RECT 449.315 3.235 449.645 3.565 ;
        RECT 449.315 1.875 449.645 2.205 ;
        RECT 449.315 0.515 449.645 0.845 ;
        RECT 449.32 -8.32 449.64 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 450.675 15.475 451.005 15.805 ;
        RECT 450.675 11.395 451.005 11.725 ;
        RECT 450.675 10.035 451.005 10.365 ;
        RECT 450.675 8.675 451.005 9.005 ;
        RECT 450.675 7.315 451.005 7.645 ;
        RECT 450.675 5.955 451.005 6.285 ;
        RECT 450.675 4.595 451.005 4.925 ;
        RECT 450.675 3.235 451.005 3.565 ;
        RECT 450.675 1.875 451.005 2.205 ;
        RECT 450.675 0.515 451.005 0.845 ;
        RECT 450.68 -8.32 451 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 452.035 15.475 452.365 15.805 ;
        RECT 452.035 10.035 452.365 10.365 ;
        RECT 452.035 8.675 452.365 9.005 ;
        RECT 452.035 7.315 452.365 7.645 ;
        RECT 452.035 5.955 452.365 6.285 ;
        RECT 452.035 4.595 452.365 4.925 ;
        RECT 452.035 3.235 452.365 3.565 ;
        RECT 452.035 1.875 452.365 2.205 ;
        RECT 452.035 0.515 452.365 0.845 ;
        RECT 452.04 -8.32 452.36 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 453.395 15.475 453.725 15.805 ;
        RECT 453.395 10.035 453.725 10.365 ;
        RECT 453.395 8.675 453.725 9.005 ;
        RECT 453.395 7.315 453.725 7.645 ;
        RECT 453.395 5.955 453.725 6.285 ;
        RECT 453.395 4.595 453.725 4.925 ;
        RECT 453.395 3.235 453.725 3.565 ;
        RECT 453.395 1.875 453.725 2.205 ;
        RECT 453.395 0.515 453.725 0.845 ;
        RECT 453.4 -8.32 453.72 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 454.755 15.475 455.085 15.805 ;
        RECT 454.755 10.035 455.085 10.365 ;
        RECT 454.755 8.675 455.085 9.005 ;
        RECT 454.755 7.315 455.085 7.645 ;
        RECT 454.755 5.955 455.085 6.285 ;
        RECT 454.755 4.595 455.085 4.925 ;
        RECT 454.755 3.235 455.085 3.565 ;
        RECT 454.755 1.875 455.085 2.205 ;
        RECT 454.755 0.515 455.085 0.845 ;
        RECT 454.76 -8.32 455.08 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 456.115 15.475 456.445 15.805 ;
        RECT 456.115 10.035 456.445 10.365 ;
        RECT 456.115 8.675 456.445 9.005 ;
        RECT 456.115 7.315 456.445 7.645 ;
        RECT 456.115 5.955 456.445 6.285 ;
        RECT 456.115 4.595 456.445 4.925 ;
        RECT 456.115 3.235 456.445 3.565 ;
        RECT 456.115 1.875 456.445 2.205 ;
        RECT 456.115 0.515 456.445 0.845 ;
        RECT 456.12 -8.32 456.44 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 457.475 15.475 457.805 15.805 ;
        RECT 457.475 10.035 457.805 10.365 ;
        RECT 457.475 8.675 457.805 9.005 ;
        RECT 457.475 7.315 457.805 7.645 ;
        RECT 457.475 5.955 457.805 6.285 ;
        RECT 457.475 4.595 457.805 4.925 ;
        RECT 457.475 3.235 457.805 3.565 ;
        RECT 457.475 1.875 457.805 2.205 ;
        RECT 457.475 0.515 457.805 0.845 ;
        RECT 457.48 -8.32 457.8 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 458.835 15.475 459.165 15.805 ;
        RECT 458.835 11.395 459.165 11.725 ;
        RECT 458.835 10.035 459.165 10.365 ;
        RECT 458.835 8.675 459.165 9.005 ;
        RECT 458.835 7.315 459.165 7.645 ;
        RECT 458.835 5.955 459.165 6.285 ;
        RECT 458.835 4.595 459.165 4.925 ;
        RECT 458.835 3.235 459.165 3.565 ;
        RECT 458.835 1.875 459.165 2.205 ;
        RECT 458.835 0.515 459.165 0.845 ;
        RECT 458.84 -8.32 459.16 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 460.195 15.475 460.525 15.805 ;
        RECT 460.195 11.395 460.525 11.725 ;
        RECT 460.195 10.035 460.525 10.365 ;
        RECT 460.195 8.675 460.525 9.005 ;
        RECT 460.195 7.315 460.525 7.645 ;
        RECT 460.195 5.955 460.525 6.285 ;
        RECT 460.195 4.595 460.525 4.925 ;
        RECT 460.195 3.235 460.525 3.565 ;
        RECT 460.195 1.875 460.525 2.205 ;
        RECT 460.195 0.515 460.525 0.845 ;
        RECT 460.2 -8.32 460.52 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 461.555 15.475 461.885 15.805 ;
        RECT 461.555 11.395 461.885 11.725 ;
        RECT 461.555 10.035 461.885 10.365 ;
        RECT 461.555 8.675 461.885 9.005 ;
        RECT 461.555 7.315 461.885 7.645 ;
        RECT 461.555 5.955 461.885 6.285 ;
        RECT 461.555 4.595 461.885 4.925 ;
        RECT 461.555 3.235 461.885 3.565 ;
        RECT 461.555 1.875 461.885 2.205 ;
        RECT 461.555 0.515 461.885 0.845 ;
        RECT 461.56 -8.32 461.88 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 462.915 15.475 463.245 15.805 ;
        RECT 462.915 10.035 463.245 10.365 ;
        RECT 462.915 8.675 463.245 9.005 ;
        RECT 462.915 7.315 463.245 7.645 ;
        RECT 462.915 5.955 463.245 6.285 ;
        RECT 462.915 4.595 463.245 4.925 ;
        RECT 462.915 3.235 463.245 3.565 ;
        RECT 462.915 1.875 463.245 2.205 ;
        RECT 462.915 0.515 463.245 0.845 ;
        RECT 462.92 -8.32 463.24 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 464.275 15.475 464.605 15.805 ;
        RECT 464.275 10.035 464.605 10.365 ;
        RECT 464.275 8.675 464.605 9.005 ;
        RECT 464.275 7.315 464.605 7.645 ;
        RECT 464.275 5.955 464.605 6.285 ;
        RECT 464.275 4.595 464.605 4.925 ;
        RECT 464.275 3.235 464.605 3.565 ;
        RECT 464.275 1.875 464.605 2.205 ;
        RECT 464.275 0.515 464.605 0.845 ;
        RECT 464.28 -8.32 464.6 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 465.635 15.475 465.965 15.805 ;
        RECT 465.635 10.035 465.965 10.365 ;
        RECT 465.635 8.675 465.965 9.005 ;
        RECT 465.635 7.315 465.965 7.645 ;
        RECT 465.635 5.955 465.965 6.285 ;
        RECT 465.635 4.595 465.965 4.925 ;
        RECT 465.635 3.235 465.965 3.565 ;
        RECT 465.635 1.875 465.965 2.205 ;
        RECT 465.635 0.515 465.965 0.845 ;
        RECT 465.64 -8.32 465.96 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 466.995 15.475 467.325 15.805 ;
        RECT 466.995 10.035 467.325 10.365 ;
        RECT 466.995 8.675 467.325 9.005 ;
        RECT 466.995 7.315 467.325 7.645 ;
        RECT 466.995 5.955 467.325 6.285 ;
        RECT 466.995 4.595 467.325 4.925 ;
        RECT 466.995 3.235 467.325 3.565 ;
        RECT 466.995 1.875 467.325 2.205 ;
        RECT 466.995 0.515 467.325 0.845 ;
        RECT 467 -8.32 467.32 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 468.355 15.475 468.685 15.805 ;
        RECT 468.355 10.035 468.685 10.365 ;
        RECT 468.355 8.675 468.685 9.005 ;
        RECT 468.355 7.315 468.685 7.645 ;
        RECT 468.355 5.955 468.685 6.285 ;
        RECT 468.355 4.595 468.685 4.925 ;
        RECT 468.355 3.235 468.685 3.565 ;
        RECT 468.355 1.875 468.685 2.205 ;
        RECT 468.355 0.515 468.685 0.845 ;
        RECT 468.36 -8.32 468.68 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 469.715 15.475 470.045 15.805 ;
        RECT 469.715 10.035 470.045 10.365 ;
        RECT 469.715 8.675 470.045 9.005 ;
        RECT 469.715 7.315 470.045 7.645 ;
        RECT 469.715 5.955 470.045 6.285 ;
        RECT 469.715 4.595 470.045 4.925 ;
        RECT 469.715 3.235 470.045 3.565 ;
        RECT 469.715 1.875 470.045 2.205 ;
        RECT 469.715 0.515 470.045 0.845 ;
        RECT 469.72 -8.32 470.04 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 471.075 15.475 471.405 15.805 ;
        RECT 471.075 11.395 471.405 11.725 ;
        RECT 471.075 10.035 471.405 10.365 ;
        RECT 471.075 8.675 471.405 9.005 ;
        RECT 471.075 7.315 471.405 7.645 ;
        RECT 471.075 5.955 471.405 6.285 ;
        RECT 471.075 4.595 471.405 4.925 ;
        RECT 471.075 3.235 471.405 3.565 ;
        RECT 471.075 1.875 471.405 2.205 ;
        RECT 471.075 0.515 471.405 0.845 ;
        RECT 471.08 -8.32 471.4 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 472.435 15.475 472.765 15.805 ;
        RECT 472.435 11.395 472.765 11.725 ;
        RECT 472.435 10.035 472.765 10.365 ;
        RECT 472.435 8.675 472.765 9.005 ;
        RECT 472.435 7.315 472.765 7.645 ;
        RECT 472.435 5.955 472.765 6.285 ;
        RECT 472.435 4.595 472.765 4.925 ;
        RECT 472.435 3.235 472.765 3.565 ;
        RECT 472.435 1.875 472.765 2.205 ;
        RECT 472.435 0.515 472.765 0.845 ;
        RECT 472.44 -8.32 472.76 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 473.795 15.475 474.125 15.805 ;
        RECT 473.795 11.395 474.125 11.725 ;
        RECT 473.795 10.035 474.125 10.365 ;
        RECT 473.795 8.675 474.125 9.005 ;
        RECT 473.795 7.315 474.125 7.645 ;
        RECT 473.795 5.955 474.125 6.285 ;
        RECT 473.795 4.595 474.125 4.925 ;
        RECT 473.795 3.235 474.125 3.565 ;
        RECT 473.795 1.875 474.125 2.205 ;
        RECT 473.795 0.515 474.125 0.845 ;
        RECT 473.8 -8.32 474.12 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 475.155 15.475 475.485 15.805 ;
        RECT 475.155 10.035 475.485 10.365 ;
        RECT 475.155 8.675 475.485 9.005 ;
        RECT 475.155 7.315 475.485 7.645 ;
        RECT 475.155 5.955 475.485 6.285 ;
        RECT 475.155 4.595 475.485 4.925 ;
        RECT 475.155 3.235 475.485 3.565 ;
        RECT 475.155 1.875 475.485 2.205 ;
        RECT 475.155 0.515 475.485 0.845 ;
        RECT 475.16 -8.32 475.48 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 476.515 15.475 476.845 15.805 ;
        RECT 476.515 10.035 476.845 10.365 ;
        RECT 476.515 8.675 476.845 9.005 ;
        RECT 476.515 7.315 476.845 7.645 ;
        RECT 476.515 5.955 476.845 6.285 ;
        RECT 476.515 4.595 476.845 4.925 ;
        RECT 476.515 3.235 476.845 3.565 ;
        RECT 476.515 1.875 476.845 2.205 ;
        RECT 476.515 0.515 476.845 0.845 ;
        RECT 476.52 -8.32 476.84 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 477.875 15.475 478.205 15.805 ;
        RECT 477.875 10.035 478.205 10.365 ;
        RECT 477.875 8.675 478.205 9.005 ;
        RECT 477.875 7.315 478.205 7.645 ;
        RECT 477.875 5.955 478.205 6.285 ;
        RECT 477.875 4.595 478.205 4.925 ;
        RECT 477.875 3.235 478.205 3.565 ;
        RECT 477.875 1.875 478.205 2.205 ;
        RECT 477.875 0.515 478.205 0.845 ;
        RECT 477.88 -8.32 478.2 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 479.235 15.475 479.565 15.805 ;
        RECT 479.235 10.035 479.565 10.365 ;
        RECT 479.235 8.675 479.565 9.005 ;
        RECT 479.235 7.315 479.565 7.645 ;
        RECT 479.235 5.955 479.565 6.285 ;
        RECT 479.235 4.595 479.565 4.925 ;
        RECT 479.235 3.235 479.565 3.565 ;
        RECT 479.235 1.875 479.565 2.205 ;
        RECT 479.235 0.515 479.565 0.845 ;
        RECT 479.24 -8.32 479.56 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 480.595 15.475 480.925 15.805 ;
        RECT 480.595 10.035 480.925 10.365 ;
        RECT 480.595 8.675 480.925 9.005 ;
        RECT 480.595 7.315 480.925 7.645 ;
        RECT 480.595 5.955 480.925 6.285 ;
        RECT 480.595 4.595 480.925 4.925 ;
        RECT 480.595 3.235 480.925 3.565 ;
        RECT 480.595 1.875 480.925 2.205 ;
        RECT 480.595 0.515 480.925 0.845 ;
        RECT 480.6 -8.32 480.92 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 481.955 15.475 482.285 15.805 ;
        RECT 481.955 10.035 482.285 10.365 ;
        RECT 481.955 8.675 482.285 9.005 ;
        RECT 481.955 7.315 482.285 7.645 ;
        RECT 481.955 5.955 482.285 6.285 ;
        RECT 481.955 4.595 482.285 4.925 ;
        RECT 481.955 3.235 482.285 3.565 ;
        RECT 481.955 1.875 482.285 2.205 ;
        RECT 481.955 0.515 482.285 0.845 ;
        RECT 481.96 -8.32 482.28 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 483.315 15.475 483.645 15.805 ;
        RECT 483.315 11.395 483.645 11.725 ;
        RECT 483.315 10.035 483.645 10.365 ;
        RECT 483.315 8.675 483.645 9.005 ;
        RECT 483.315 7.315 483.645 7.645 ;
        RECT 483.315 5.955 483.645 6.285 ;
        RECT 483.315 4.595 483.645 4.925 ;
        RECT 483.315 3.235 483.645 3.565 ;
        RECT 483.315 1.875 483.645 2.205 ;
        RECT 483.315 0.515 483.645 0.845 ;
        RECT 483.32 -8.32 483.64 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 484.675 15.475 485.005 15.805 ;
        RECT 484.675 11.395 485.005 11.725 ;
        RECT 484.675 10.035 485.005 10.365 ;
        RECT 484.675 8.675 485.005 9.005 ;
        RECT 484.675 7.315 485.005 7.645 ;
        RECT 484.675 5.955 485.005 6.285 ;
        RECT 484.675 4.595 485.005 4.925 ;
        RECT 484.675 3.235 485.005 3.565 ;
        RECT 484.675 1.875 485.005 2.205 ;
        RECT 484.675 0.515 485.005 0.845 ;
        RECT 484.68 -8.32 485 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 486.035 15.475 486.365 15.805 ;
        RECT 486.035 11.395 486.365 11.725 ;
        RECT 486.035 10.035 486.365 10.365 ;
        RECT 486.035 8.675 486.365 9.005 ;
        RECT 486.035 7.315 486.365 7.645 ;
        RECT 486.035 5.955 486.365 6.285 ;
        RECT 486.035 4.595 486.365 4.925 ;
        RECT 486.035 3.235 486.365 3.565 ;
        RECT 486.035 1.875 486.365 2.205 ;
        RECT 486.035 0.515 486.365 0.845 ;
        RECT 486.04 -8.32 486.36 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 487.395 15.475 487.725 15.805 ;
        RECT 487.395 10.035 487.725 10.365 ;
        RECT 487.395 8.675 487.725 9.005 ;
        RECT 487.395 7.315 487.725 7.645 ;
        RECT 487.395 5.955 487.725 6.285 ;
        RECT 487.395 4.595 487.725 4.925 ;
        RECT 487.395 3.235 487.725 3.565 ;
        RECT 487.395 1.875 487.725 2.205 ;
        RECT 487.395 0.515 487.725 0.845 ;
        RECT 487.4 -8.32 487.72 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 488.755 15.475 489.085 15.805 ;
        RECT 488.755 10.035 489.085 10.365 ;
        RECT 488.755 8.675 489.085 9.005 ;
        RECT 488.755 7.315 489.085 7.645 ;
        RECT 488.755 5.955 489.085 6.285 ;
        RECT 488.755 4.595 489.085 4.925 ;
        RECT 488.755 3.235 489.085 3.565 ;
        RECT 488.755 1.875 489.085 2.205 ;
        RECT 488.755 0.515 489.085 0.845 ;
        RECT 488.76 -8.32 489.08 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 490.115 15.475 490.445 15.805 ;
        RECT 490.115 10.035 490.445 10.365 ;
        RECT 490.115 8.675 490.445 9.005 ;
        RECT 490.115 7.315 490.445 7.645 ;
        RECT 490.115 5.955 490.445 6.285 ;
        RECT 490.115 4.595 490.445 4.925 ;
        RECT 490.115 3.235 490.445 3.565 ;
        RECT 490.115 1.875 490.445 2.205 ;
        RECT 490.115 0.515 490.445 0.845 ;
        RECT 490.12 -8.32 490.44 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 491.475 15.475 491.805 15.805 ;
        RECT 491.475 10.035 491.805 10.365 ;
        RECT 491.475 8.675 491.805 9.005 ;
        RECT 491.475 7.315 491.805 7.645 ;
        RECT 491.475 5.955 491.805 6.285 ;
        RECT 491.475 4.595 491.805 4.925 ;
        RECT 491.475 3.235 491.805 3.565 ;
        RECT 491.475 1.875 491.805 2.205 ;
        RECT 491.475 0.515 491.805 0.845 ;
        RECT 491.48 -8.32 491.8 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 492.835 15.475 493.165 15.805 ;
        RECT 492.835 10.035 493.165 10.365 ;
        RECT 492.835 8.675 493.165 9.005 ;
        RECT 492.835 7.315 493.165 7.645 ;
        RECT 492.835 5.955 493.165 6.285 ;
        RECT 492.835 4.595 493.165 4.925 ;
        RECT 492.835 3.235 493.165 3.565 ;
        RECT 492.835 1.875 493.165 2.205 ;
        RECT 492.835 0.515 493.165 0.845 ;
        RECT 492.84 -8.32 493.16 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 494.195 15.475 494.525 15.805 ;
        RECT 494.195 10.035 494.525 10.365 ;
        RECT 494.195 8.675 494.525 9.005 ;
        RECT 494.195 7.315 494.525 7.645 ;
        RECT 494.195 5.955 494.525 6.285 ;
        RECT 494.195 4.595 494.525 4.925 ;
        RECT 494.195 3.235 494.525 3.565 ;
        RECT 494.195 1.875 494.525 2.205 ;
        RECT 494.195 0.515 494.525 0.845 ;
        RECT 494.2 -8.32 494.52 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 495.555 15.475 495.885 15.805 ;
        RECT 495.555 11.395 495.885 11.725 ;
        RECT 495.555 10.035 495.885 10.365 ;
        RECT 495.555 8.675 495.885 9.005 ;
        RECT 495.555 7.315 495.885 7.645 ;
        RECT 495.555 5.955 495.885 6.285 ;
        RECT 495.555 4.595 495.885 4.925 ;
        RECT 495.555 3.235 495.885 3.565 ;
        RECT 495.555 1.875 495.885 2.205 ;
        RECT 495.555 0.515 495.885 0.845 ;
        RECT 495.56 -8.32 495.88 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 496.915 15.475 497.245 15.805 ;
        RECT 496.915 11.395 497.245 11.725 ;
        RECT 496.915 10.035 497.245 10.365 ;
        RECT 496.915 8.675 497.245 9.005 ;
        RECT 496.915 7.315 497.245 7.645 ;
        RECT 496.915 5.955 497.245 6.285 ;
        RECT 496.915 4.595 497.245 4.925 ;
        RECT 496.915 3.235 497.245 3.565 ;
        RECT 496.915 1.875 497.245 2.205 ;
        RECT 496.915 0.515 497.245 0.845 ;
        RECT 496.92 -8.32 497.24 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 498.275 15.475 498.605 15.805 ;
        RECT 498.275 11.395 498.605 11.725 ;
        RECT 498.275 10.035 498.605 10.365 ;
        RECT 498.275 8.675 498.605 9.005 ;
        RECT 498.275 7.315 498.605 7.645 ;
        RECT 498.275 5.955 498.605 6.285 ;
        RECT 498.275 4.595 498.605 4.925 ;
        RECT 498.275 3.235 498.605 3.565 ;
        RECT 498.275 1.875 498.605 2.205 ;
        RECT 498.275 0.515 498.605 0.845 ;
        RECT 498.28 -8.32 498.6 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 499.635 15.475 499.965 15.805 ;
        RECT 499.635 10.035 499.965 10.365 ;
        RECT 499.635 8.675 499.965 9.005 ;
        RECT 499.635 7.315 499.965 7.645 ;
        RECT 499.635 5.955 499.965 6.285 ;
        RECT 499.635 4.595 499.965 4.925 ;
        RECT 499.635 3.235 499.965 3.565 ;
        RECT 499.635 1.875 499.965 2.205 ;
        RECT 499.635 0.515 499.965 0.845 ;
        RECT 499.64 -8.32 499.96 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 500.995 15.475 501.325 15.805 ;
        RECT 500.995 10.035 501.325 10.365 ;
        RECT 500.995 8.675 501.325 9.005 ;
        RECT 500.995 7.315 501.325 7.645 ;
        RECT 500.995 5.955 501.325 6.285 ;
        RECT 500.995 4.595 501.325 4.925 ;
        RECT 500.995 3.235 501.325 3.565 ;
        RECT 500.995 1.875 501.325 2.205 ;
        RECT 500.995 0.515 501.325 0.845 ;
        RECT 501 -8.32 501.32 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 502.355 15.475 502.685 15.805 ;
        RECT 502.355 10.035 502.685 10.365 ;
        RECT 502.355 8.675 502.685 9.005 ;
        RECT 502.355 7.315 502.685 7.645 ;
        RECT 502.355 5.955 502.685 6.285 ;
        RECT 502.355 4.595 502.685 4.925 ;
        RECT 502.355 3.235 502.685 3.565 ;
        RECT 502.355 1.875 502.685 2.205 ;
        RECT 502.355 0.515 502.685 0.845 ;
        RECT 502.36 -8.32 502.68 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 503.715 15.475 504.045 15.805 ;
        RECT 503.715 10.035 504.045 10.365 ;
        RECT 503.715 8.675 504.045 9.005 ;
        RECT 503.715 7.315 504.045 7.645 ;
        RECT 503.715 5.955 504.045 6.285 ;
        RECT 503.715 4.595 504.045 4.925 ;
        RECT 503.715 3.235 504.045 3.565 ;
        RECT 503.715 1.875 504.045 2.205 ;
        RECT 503.715 0.515 504.045 0.845 ;
        RECT 503.72 -8.32 504.04 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 505.075 15.475 505.405 15.805 ;
        RECT 505.075 10.035 505.405 10.365 ;
        RECT 505.075 8.675 505.405 9.005 ;
        RECT 505.075 7.315 505.405 7.645 ;
        RECT 505.075 5.955 505.405 6.285 ;
        RECT 505.075 4.595 505.405 4.925 ;
        RECT 505.075 3.235 505.405 3.565 ;
        RECT 505.075 1.875 505.405 2.205 ;
        RECT 505.075 0.515 505.405 0.845 ;
        RECT 505.08 -8.32 505.4 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 506.435 15.475 506.765 15.805 ;
        RECT 506.435 10.035 506.765 10.365 ;
        RECT 506.435 8.675 506.765 9.005 ;
        RECT 506.435 7.315 506.765 7.645 ;
        RECT 506.435 5.955 506.765 6.285 ;
        RECT 506.435 4.595 506.765 4.925 ;
        RECT 506.435 3.235 506.765 3.565 ;
        RECT 506.435 1.875 506.765 2.205 ;
        RECT 506.435 0.515 506.765 0.845 ;
        RECT 506.44 -8.32 506.76 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 507.795 7.315 508.125 7.645 ;
        RECT 507.795 5.955 508.125 6.285 ;
        RECT 507.795 4.595 508.125 4.925 ;
        RECT 507.795 3.235 508.125 3.565 ;
        RECT 507.795 1.875 508.125 2.205 ;
        RECT 507.795 0.515 508.125 0.845 ;
        RECT 507.8 -8.32 508.12 15.805 ;
        RECT 507.795 15.475 508.125 15.805 ;
        RECT 507.795 11.395 508.125 11.725 ;
        RECT 507.795 10.035 508.125 10.365 ;
        RECT 507.795 8.675 508.125 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 246.675 15.475 247.005 15.805 ;
        RECT 246.675 11.395 247.005 11.725 ;
        RECT 246.675 10.035 247.005 10.365 ;
        RECT 246.675 8.675 247.005 9.005 ;
        RECT 246.675 7.315 247.005 7.645 ;
        RECT 246.675 5.955 247.005 6.285 ;
        RECT 246.675 4.595 247.005 4.925 ;
        RECT 246.675 3.235 247.005 3.565 ;
        RECT 246.675 1.875 247.005 2.205 ;
        RECT 246.675 0.515 247.005 0.845 ;
        RECT 246.68 -8.32 247 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.035 15.475 248.365 15.805 ;
        RECT 248.035 10.035 248.365 10.365 ;
        RECT 248.035 8.675 248.365 9.005 ;
        RECT 248.035 7.315 248.365 7.645 ;
        RECT 248.035 5.955 248.365 6.285 ;
        RECT 248.035 4.595 248.365 4.925 ;
        RECT 248.035 3.235 248.365 3.565 ;
        RECT 248.035 1.875 248.365 2.205 ;
        RECT 248.035 0.515 248.365 0.845 ;
        RECT 248.04 -8.32 248.36 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 249.395 15.475 249.725 15.805 ;
        RECT 249.395 10.035 249.725 10.365 ;
        RECT 249.395 8.675 249.725 9.005 ;
        RECT 249.395 7.315 249.725 7.645 ;
        RECT 249.395 5.955 249.725 6.285 ;
        RECT 249.395 4.595 249.725 4.925 ;
        RECT 249.395 3.235 249.725 3.565 ;
        RECT 249.395 1.875 249.725 2.205 ;
        RECT 249.395 0.515 249.725 0.845 ;
        RECT 249.4 -8.32 249.72 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.755 15.475 251.085 15.805 ;
        RECT 250.755 10.035 251.085 10.365 ;
        RECT 250.755 8.675 251.085 9.005 ;
        RECT 250.755 7.315 251.085 7.645 ;
        RECT 250.755 5.955 251.085 6.285 ;
        RECT 250.755 4.595 251.085 4.925 ;
        RECT 250.755 3.235 251.085 3.565 ;
        RECT 250.755 1.875 251.085 2.205 ;
        RECT 250.755 0.515 251.085 0.845 ;
        RECT 250.76 -8.32 251.08 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.115 15.475 252.445 15.805 ;
        RECT 252.115 10.035 252.445 10.365 ;
        RECT 252.115 8.675 252.445 9.005 ;
        RECT 252.115 7.315 252.445 7.645 ;
        RECT 252.115 5.955 252.445 6.285 ;
        RECT 252.115 4.595 252.445 4.925 ;
        RECT 252.115 3.235 252.445 3.565 ;
        RECT 252.115 1.875 252.445 2.205 ;
        RECT 252.115 0.515 252.445 0.845 ;
        RECT 252.12 -8.32 252.44 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 253.475 15.475 253.805 15.805 ;
        RECT 253.475 10.035 253.805 10.365 ;
        RECT 253.475 8.675 253.805 9.005 ;
        RECT 253.475 7.315 253.805 7.645 ;
        RECT 253.475 5.955 253.805 6.285 ;
        RECT 253.475 4.595 253.805 4.925 ;
        RECT 253.475 3.235 253.805 3.565 ;
        RECT 253.475 1.875 253.805 2.205 ;
        RECT 253.475 0.515 253.805 0.845 ;
        RECT 253.48 -8.32 253.8 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 254.835 15.475 255.165 15.805 ;
        RECT 254.835 11.395 255.165 11.725 ;
        RECT 254.835 10.035 255.165 10.365 ;
        RECT 254.835 8.675 255.165 9.005 ;
        RECT 254.835 7.315 255.165 7.645 ;
        RECT 254.835 5.955 255.165 6.285 ;
        RECT 254.835 4.595 255.165 4.925 ;
        RECT 254.835 3.235 255.165 3.565 ;
        RECT 254.835 1.875 255.165 2.205 ;
        RECT 254.835 0.515 255.165 0.845 ;
        RECT 254.84 -8.32 255.16 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 256.195 15.475 256.525 15.805 ;
        RECT 256.195 11.395 256.525 11.725 ;
        RECT 256.195 10.035 256.525 10.365 ;
        RECT 256.195 8.675 256.525 9.005 ;
        RECT 256.195 7.315 256.525 7.645 ;
        RECT 256.195 5.955 256.525 6.285 ;
        RECT 256.195 4.595 256.525 4.925 ;
        RECT 256.195 3.235 256.525 3.565 ;
        RECT 256.195 1.875 256.525 2.205 ;
        RECT 256.195 0.515 256.525 0.845 ;
        RECT 256.2 -8.32 256.52 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 257.555 15.475 257.885 15.805 ;
        RECT 257.555 11.395 257.885 11.725 ;
        RECT 257.555 10.035 257.885 10.365 ;
        RECT 257.555 8.675 257.885 9.005 ;
        RECT 257.555 7.315 257.885 7.645 ;
        RECT 257.555 5.955 257.885 6.285 ;
        RECT 257.555 4.595 257.885 4.925 ;
        RECT 257.555 3.235 257.885 3.565 ;
        RECT 257.555 1.875 257.885 2.205 ;
        RECT 257.555 0.515 257.885 0.845 ;
        RECT 257.56 -8.32 257.88 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.915 15.475 259.245 15.805 ;
        RECT 258.915 10.035 259.245 10.365 ;
        RECT 258.915 8.675 259.245 9.005 ;
        RECT 258.915 7.315 259.245 7.645 ;
        RECT 258.915 5.955 259.245 6.285 ;
        RECT 258.915 4.595 259.245 4.925 ;
        RECT 258.915 3.235 259.245 3.565 ;
        RECT 258.915 1.875 259.245 2.205 ;
        RECT 258.915 0.515 259.245 0.845 ;
        RECT 258.92 -8.32 259.24 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.275 15.475 260.605 15.805 ;
        RECT 260.275 10.035 260.605 10.365 ;
        RECT 260.275 8.675 260.605 9.005 ;
        RECT 260.275 7.315 260.605 7.645 ;
        RECT 260.275 5.955 260.605 6.285 ;
        RECT 260.275 4.595 260.605 4.925 ;
        RECT 260.275 3.235 260.605 3.565 ;
        RECT 260.275 1.875 260.605 2.205 ;
        RECT 260.275 0.515 260.605 0.845 ;
        RECT 260.28 -8.32 260.6 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 261.635 15.475 261.965 15.805 ;
        RECT 261.635 10.035 261.965 10.365 ;
        RECT 261.635 8.675 261.965 9.005 ;
        RECT 261.635 7.315 261.965 7.645 ;
        RECT 261.635 5.955 261.965 6.285 ;
        RECT 261.635 4.595 261.965 4.925 ;
        RECT 261.635 3.235 261.965 3.565 ;
        RECT 261.635 1.875 261.965 2.205 ;
        RECT 261.635 0.515 261.965 0.845 ;
        RECT 261.64 -8.32 261.96 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.995 15.475 263.325 15.805 ;
        RECT 262.995 10.035 263.325 10.365 ;
        RECT 262.995 8.675 263.325 9.005 ;
        RECT 262.995 7.315 263.325 7.645 ;
        RECT 262.995 5.955 263.325 6.285 ;
        RECT 262.995 4.595 263.325 4.925 ;
        RECT 262.995 3.235 263.325 3.565 ;
        RECT 262.995 1.875 263.325 2.205 ;
        RECT 262.995 0.515 263.325 0.845 ;
        RECT 263 -8.32 263.32 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 264.355 15.475 264.685 15.805 ;
        RECT 264.355 10.035 264.685 10.365 ;
        RECT 264.355 8.675 264.685 9.005 ;
        RECT 264.355 7.315 264.685 7.645 ;
        RECT 264.355 5.955 264.685 6.285 ;
        RECT 264.355 4.595 264.685 4.925 ;
        RECT 264.355 3.235 264.685 3.565 ;
        RECT 264.355 1.875 264.685 2.205 ;
        RECT 264.355 0.515 264.685 0.845 ;
        RECT 264.36 -8.32 264.68 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 265.715 15.475 266.045 15.805 ;
        RECT 265.715 10.035 266.045 10.365 ;
        RECT 265.715 8.675 266.045 9.005 ;
        RECT 265.715 7.315 266.045 7.645 ;
        RECT 265.715 5.955 266.045 6.285 ;
        RECT 265.715 4.595 266.045 4.925 ;
        RECT 265.715 3.235 266.045 3.565 ;
        RECT 265.715 1.875 266.045 2.205 ;
        RECT 265.715 0.515 266.045 0.845 ;
        RECT 265.72 -8.32 266.04 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 267.075 15.475 267.405 15.805 ;
        RECT 267.075 11.395 267.405 11.725 ;
        RECT 267.075 10.035 267.405 10.365 ;
        RECT 267.075 8.675 267.405 9.005 ;
        RECT 267.075 7.315 267.405 7.645 ;
        RECT 267.075 5.955 267.405 6.285 ;
        RECT 267.075 4.595 267.405 4.925 ;
        RECT 267.075 3.235 267.405 3.565 ;
        RECT 267.075 1.875 267.405 2.205 ;
        RECT 267.075 0.515 267.405 0.845 ;
        RECT 267.08 -8.32 267.4 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 268.435 15.475 268.765 15.805 ;
        RECT 268.435 11.395 268.765 11.725 ;
        RECT 268.435 10.035 268.765 10.365 ;
        RECT 268.435 8.675 268.765 9.005 ;
        RECT 268.435 7.315 268.765 7.645 ;
        RECT 268.435 5.955 268.765 6.285 ;
        RECT 268.435 4.595 268.765 4.925 ;
        RECT 268.435 3.235 268.765 3.565 ;
        RECT 268.435 1.875 268.765 2.205 ;
        RECT 268.435 0.515 268.765 0.845 ;
        RECT 268.44 -8.32 268.76 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.795 15.475 270.125 15.805 ;
        RECT 269.795 11.395 270.125 11.725 ;
        RECT 269.795 10.035 270.125 10.365 ;
        RECT 269.795 8.675 270.125 9.005 ;
        RECT 269.795 7.315 270.125 7.645 ;
        RECT 269.795 5.955 270.125 6.285 ;
        RECT 269.795 4.595 270.125 4.925 ;
        RECT 269.795 3.235 270.125 3.565 ;
        RECT 269.795 1.875 270.125 2.205 ;
        RECT 269.795 0.515 270.125 0.845 ;
        RECT 269.8 -8.32 270.12 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.155 15.475 271.485 15.805 ;
        RECT 271.155 10.035 271.485 10.365 ;
        RECT 271.155 8.675 271.485 9.005 ;
        RECT 271.155 7.315 271.485 7.645 ;
        RECT 271.155 5.955 271.485 6.285 ;
        RECT 271.155 4.595 271.485 4.925 ;
        RECT 271.155 3.235 271.485 3.565 ;
        RECT 271.155 1.875 271.485 2.205 ;
        RECT 271.155 0.515 271.485 0.845 ;
        RECT 271.16 -8.32 271.48 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 272.515 15.475 272.845 15.805 ;
        RECT 272.515 10.035 272.845 10.365 ;
        RECT 272.515 8.675 272.845 9.005 ;
        RECT 272.515 7.315 272.845 7.645 ;
        RECT 272.515 5.955 272.845 6.285 ;
        RECT 272.515 4.595 272.845 4.925 ;
        RECT 272.515 3.235 272.845 3.565 ;
        RECT 272.515 1.875 272.845 2.205 ;
        RECT 272.515 0.515 272.845 0.845 ;
        RECT 272.52 -8.32 272.84 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.875 15.475 274.205 15.805 ;
        RECT 273.875 10.035 274.205 10.365 ;
        RECT 273.875 8.675 274.205 9.005 ;
        RECT 273.875 7.315 274.205 7.645 ;
        RECT 273.875 5.955 274.205 6.285 ;
        RECT 273.875 4.595 274.205 4.925 ;
        RECT 273.875 3.235 274.205 3.565 ;
        RECT 273.875 1.875 274.205 2.205 ;
        RECT 273.875 0.515 274.205 0.845 ;
        RECT 273.88 -8.32 274.2 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.235 15.475 275.565 15.805 ;
        RECT 275.235 10.035 275.565 10.365 ;
        RECT 275.235 8.675 275.565 9.005 ;
        RECT 275.235 7.315 275.565 7.645 ;
        RECT 275.235 5.955 275.565 6.285 ;
        RECT 275.235 4.595 275.565 4.925 ;
        RECT 275.235 3.235 275.565 3.565 ;
        RECT 275.235 1.875 275.565 2.205 ;
        RECT 275.235 0.515 275.565 0.845 ;
        RECT 275.24 -8.32 275.56 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 276.595 15.475 276.925 15.805 ;
        RECT 276.595 10.035 276.925 10.365 ;
        RECT 276.595 8.675 276.925 9.005 ;
        RECT 276.595 7.315 276.925 7.645 ;
        RECT 276.595 5.955 276.925 6.285 ;
        RECT 276.595 4.595 276.925 4.925 ;
        RECT 276.595 3.235 276.925 3.565 ;
        RECT 276.595 1.875 276.925 2.205 ;
        RECT 276.595 0.515 276.925 0.845 ;
        RECT 276.6 -8.32 276.92 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 277.955 15.475 278.285 15.805 ;
        RECT 277.955 10.035 278.285 10.365 ;
        RECT 277.955 8.675 278.285 9.005 ;
        RECT 277.955 7.315 278.285 7.645 ;
        RECT 277.955 5.955 278.285 6.285 ;
        RECT 277.955 4.595 278.285 4.925 ;
        RECT 277.955 3.235 278.285 3.565 ;
        RECT 277.955 1.875 278.285 2.205 ;
        RECT 277.955 0.515 278.285 0.845 ;
        RECT 277.96 -8.32 278.28 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.315 15.475 279.645 15.805 ;
        RECT 279.315 11.395 279.645 11.725 ;
        RECT 279.315 10.035 279.645 10.365 ;
        RECT 279.315 8.675 279.645 9.005 ;
        RECT 279.315 7.315 279.645 7.645 ;
        RECT 279.315 5.955 279.645 6.285 ;
        RECT 279.315 4.595 279.645 4.925 ;
        RECT 279.315 3.235 279.645 3.565 ;
        RECT 279.315 1.875 279.645 2.205 ;
        RECT 279.315 0.515 279.645 0.845 ;
        RECT 279.32 -8.32 279.64 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 280.675 15.475 281.005 15.805 ;
        RECT 280.675 11.395 281.005 11.725 ;
        RECT 280.675 10.035 281.005 10.365 ;
        RECT 280.675 8.675 281.005 9.005 ;
        RECT 280.675 7.315 281.005 7.645 ;
        RECT 280.675 5.955 281.005 6.285 ;
        RECT 280.675 4.595 281.005 4.925 ;
        RECT 280.675 3.235 281.005 3.565 ;
        RECT 280.675 1.875 281.005 2.205 ;
        RECT 280.675 0.515 281.005 0.845 ;
        RECT 280.68 -8.32 281 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.035 15.475 282.365 15.805 ;
        RECT 282.035 11.395 282.365 11.725 ;
        RECT 282.035 10.035 282.365 10.365 ;
        RECT 282.035 8.675 282.365 9.005 ;
        RECT 282.035 7.315 282.365 7.645 ;
        RECT 282.035 5.955 282.365 6.285 ;
        RECT 282.035 4.595 282.365 4.925 ;
        RECT 282.035 3.235 282.365 3.565 ;
        RECT 282.035 1.875 282.365 2.205 ;
        RECT 282.035 0.515 282.365 0.845 ;
        RECT 282.04 -8.32 282.36 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 283.395 15.475 283.725 15.805 ;
        RECT 283.395 10.035 283.725 10.365 ;
        RECT 283.395 8.675 283.725 9.005 ;
        RECT 283.395 7.315 283.725 7.645 ;
        RECT 283.395 5.955 283.725 6.285 ;
        RECT 283.395 4.595 283.725 4.925 ;
        RECT 283.395 3.235 283.725 3.565 ;
        RECT 283.395 1.875 283.725 2.205 ;
        RECT 283.395 0.515 283.725 0.845 ;
        RECT 283.4 -8.32 283.72 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 284.755 15.475 285.085 15.805 ;
        RECT 284.755 10.035 285.085 10.365 ;
        RECT 284.755 8.675 285.085 9.005 ;
        RECT 284.755 7.315 285.085 7.645 ;
        RECT 284.755 5.955 285.085 6.285 ;
        RECT 284.755 4.595 285.085 4.925 ;
        RECT 284.755 3.235 285.085 3.565 ;
        RECT 284.755 1.875 285.085 2.205 ;
        RECT 284.755 0.515 285.085 0.845 ;
        RECT 284.76 -8.32 285.08 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.115 15.475 286.445 15.805 ;
        RECT 286.115 10.035 286.445 10.365 ;
        RECT 286.115 8.675 286.445 9.005 ;
        RECT 286.115 7.315 286.445 7.645 ;
        RECT 286.115 5.955 286.445 6.285 ;
        RECT 286.115 4.595 286.445 4.925 ;
        RECT 286.115 3.235 286.445 3.565 ;
        RECT 286.115 1.875 286.445 2.205 ;
        RECT 286.115 0.515 286.445 0.845 ;
        RECT 286.12 -8.32 286.44 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 287.475 15.475 287.805 15.805 ;
        RECT 287.475 10.035 287.805 10.365 ;
        RECT 287.475 8.675 287.805 9.005 ;
        RECT 287.475 7.315 287.805 7.645 ;
        RECT 287.475 5.955 287.805 6.285 ;
        RECT 287.475 4.595 287.805 4.925 ;
        RECT 287.475 3.235 287.805 3.565 ;
        RECT 287.475 1.875 287.805 2.205 ;
        RECT 287.475 0.515 287.805 0.845 ;
        RECT 287.48 -8.32 287.8 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.835 15.475 289.165 15.805 ;
        RECT 288.835 10.035 289.165 10.365 ;
        RECT 288.835 8.675 289.165 9.005 ;
        RECT 288.835 7.315 289.165 7.645 ;
        RECT 288.835 5.955 289.165 6.285 ;
        RECT 288.835 4.595 289.165 4.925 ;
        RECT 288.835 3.235 289.165 3.565 ;
        RECT 288.835 1.875 289.165 2.205 ;
        RECT 288.835 0.515 289.165 0.845 ;
        RECT 288.84 -8.32 289.16 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.195 15.475 290.525 15.805 ;
        RECT 290.195 10.035 290.525 10.365 ;
        RECT 290.195 8.675 290.525 9.005 ;
        RECT 290.195 7.315 290.525 7.645 ;
        RECT 290.195 5.955 290.525 6.285 ;
        RECT 290.195 4.595 290.525 4.925 ;
        RECT 290.195 3.235 290.525 3.565 ;
        RECT 290.195 1.875 290.525 2.205 ;
        RECT 290.195 0.515 290.525 0.845 ;
        RECT 290.2 -8.32 290.52 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 291.555 15.475 291.885 15.805 ;
        RECT 291.555 11.395 291.885 11.725 ;
        RECT 291.555 10.035 291.885 10.365 ;
        RECT 291.555 8.675 291.885 9.005 ;
        RECT 291.555 7.315 291.885 7.645 ;
        RECT 291.555 5.955 291.885 6.285 ;
        RECT 291.555 4.595 291.885 4.925 ;
        RECT 291.555 3.235 291.885 3.565 ;
        RECT 291.555 1.875 291.885 2.205 ;
        RECT 291.555 0.515 291.885 0.845 ;
        RECT 291.56 -8.32 291.88 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.915 15.475 293.245 15.805 ;
        RECT 292.915 11.395 293.245 11.725 ;
        RECT 292.915 10.035 293.245 10.365 ;
        RECT 292.915 8.675 293.245 9.005 ;
        RECT 292.915 7.315 293.245 7.645 ;
        RECT 292.915 5.955 293.245 6.285 ;
        RECT 292.915 4.595 293.245 4.925 ;
        RECT 292.915 3.235 293.245 3.565 ;
        RECT 292.915 1.875 293.245 2.205 ;
        RECT 292.915 0.515 293.245 0.845 ;
        RECT 292.92 -8.32 293.24 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.275 15.475 294.605 15.805 ;
        RECT 294.275 11.395 294.605 11.725 ;
        RECT 294.275 10.035 294.605 10.365 ;
        RECT 294.275 8.675 294.605 9.005 ;
        RECT 294.275 7.315 294.605 7.645 ;
        RECT 294.275 5.955 294.605 6.285 ;
        RECT 294.275 4.595 294.605 4.925 ;
        RECT 294.275 3.235 294.605 3.565 ;
        RECT 294.275 1.875 294.605 2.205 ;
        RECT 294.275 0.515 294.605 0.845 ;
        RECT 294.28 -8.32 294.6 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 295.635 15.475 295.965 15.805 ;
        RECT 295.635 10.035 295.965 10.365 ;
        RECT 295.635 8.675 295.965 9.005 ;
        RECT 295.635 7.315 295.965 7.645 ;
        RECT 295.635 5.955 295.965 6.285 ;
        RECT 295.635 4.595 295.965 4.925 ;
        RECT 295.635 3.235 295.965 3.565 ;
        RECT 295.635 1.875 295.965 2.205 ;
        RECT 295.635 0.515 295.965 0.845 ;
        RECT 295.64 -8.32 295.96 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 296.995 15.475 297.325 15.805 ;
        RECT 296.995 10.035 297.325 10.365 ;
        RECT 296.995 8.675 297.325 9.005 ;
        RECT 296.995 7.315 297.325 7.645 ;
        RECT 296.995 5.955 297.325 6.285 ;
        RECT 296.995 4.595 297.325 4.925 ;
        RECT 296.995 3.235 297.325 3.565 ;
        RECT 296.995 1.875 297.325 2.205 ;
        RECT 296.995 0.515 297.325 0.845 ;
        RECT 297 -8.32 297.32 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 298.355 15.475 298.685 15.805 ;
        RECT 298.355 10.035 298.685 10.365 ;
        RECT 298.355 8.675 298.685 9.005 ;
        RECT 298.355 7.315 298.685 7.645 ;
        RECT 298.355 5.955 298.685 6.285 ;
        RECT 298.355 4.595 298.685 4.925 ;
        RECT 298.355 3.235 298.685 3.565 ;
        RECT 298.355 1.875 298.685 2.205 ;
        RECT 298.355 0.515 298.685 0.845 ;
        RECT 298.36 -8.32 298.68 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 299.715 15.475 300.045 15.805 ;
        RECT 299.715 10.035 300.045 10.365 ;
        RECT 299.715 8.675 300.045 9.005 ;
        RECT 299.715 7.315 300.045 7.645 ;
        RECT 299.715 5.955 300.045 6.285 ;
        RECT 299.715 4.595 300.045 4.925 ;
        RECT 299.715 3.235 300.045 3.565 ;
        RECT 299.715 1.875 300.045 2.205 ;
        RECT 299.715 0.515 300.045 0.845 ;
        RECT 299.72 -8.32 300.04 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.075 15.475 301.405 15.805 ;
        RECT 301.075 10.035 301.405 10.365 ;
        RECT 301.075 8.675 301.405 9.005 ;
        RECT 301.075 7.315 301.405 7.645 ;
        RECT 301.075 5.955 301.405 6.285 ;
        RECT 301.075 4.595 301.405 4.925 ;
        RECT 301.075 3.235 301.405 3.565 ;
        RECT 301.075 1.875 301.405 2.205 ;
        RECT 301.075 0.515 301.405 0.845 ;
        RECT 301.08 -8.32 301.4 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 302.435 15.475 302.765 15.805 ;
        RECT 302.435 10.035 302.765 10.365 ;
        RECT 302.435 8.675 302.765 9.005 ;
        RECT 302.435 7.315 302.765 7.645 ;
        RECT 302.435 5.955 302.765 6.285 ;
        RECT 302.435 4.595 302.765 4.925 ;
        RECT 302.435 3.235 302.765 3.565 ;
        RECT 302.435 1.875 302.765 2.205 ;
        RECT 302.435 0.515 302.765 0.845 ;
        RECT 302.44 -8.32 302.76 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.795 15.475 304.125 15.805 ;
        RECT 303.795 11.395 304.125 11.725 ;
        RECT 303.795 10.035 304.125 10.365 ;
        RECT 303.795 8.675 304.125 9.005 ;
        RECT 303.795 7.315 304.125 7.645 ;
        RECT 303.795 5.955 304.125 6.285 ;
        RECT 303.795 4.595 304.125 4.925 ;
        RECT 303.795 3.235 304.125 3.565 ;
        RECT 303.795 1.875 304.125 2.205 ;
        RECT 303.795 0.515 304.125 0.845 ;
        RECT 303.8 -8.32 304.12 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.155 15.475 305.485 15.805 ;
        RECT 305.155 11.395 305.485 11.725 ;
        RECT 305.155 10.035 305.485 10.365 ;
        RECT 305.155 8.675 305.485 9.005 ;
        RECT 305.155 7.315 305.485 7.645 ;
        RECT 305.155 5.955 305.485 6.285 ;
        RECT 305.155 4.595 305.485 4.925 ;
        RECT 305.155 3.235 305.485 3.565 ;
        RECT 305.155 1.875 305.485 2.205 ;
        RECT 305.155 0.515 305.485 0.845 ;
        RECT 305.16 -8.32 305.48 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 306.515 15.475 306.845 15.805 ;
        RECT 306.515 11.395 306.845 11.725 ;
        RECT 306.515 10.035 306.845 10.365 ;
        RECT 306.515 8.675 306.845 9.005 ;
        RECT 306.515 7.315 306.845 7.645 ;
        RECT 306.515 5.955 306.845 6.285 ;
        RECT 306.515 4.595 306.845 4.925 ;
        RECT 306.515 3.235 306.845 3.565 ;
        RECT 306.515 1.875 306.845 2.205 ;
        RECT 306.515 0.515 306.845 0.845 ;
        RECT 306.52 -8.32 306.84 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.875 15.475 308.205 15.805 ;
        RECT 307.875 10.035 308.205 10.365 ;
        RECT 307.875 8.675 308.205 9.005 ;
        RECT 307.875 7.315 308.205 7.645 ;
        RECT 307.875 5.955 308.205 6.285 ;
        RECT 307.875 4.595 308.205 4.925 ;
        RECT 307.875 3.235 308.205 3.565 ;
        RECT 307.875 1.875 308.205 2.205 ;
        RECT 307.875 0.515 308.205 0.845 ;
        RECT 307.88 -8.32 308.2 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.235 15.475 309.565 15.805 ;
        RECT 309.235 10.035 309.565 10.365 ;
        RECT 309.235 8.675 309.565 9.005 ;
        RECT 309.235 7.315 309.565 7.645 ;
        RECT 309.235 5.955 309.565 6.285 ;
        RECT 309.235 4.595 309.565 4.925 ;
        RECT 309.235 3.235 309.565 3.565 ;
        RECT 309.235 1.875 309.565 2.205 ;
        RECT 309.235 0.515 309.565 0.845 ;
        RECT 309.24 -8.32 309.56 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 310.595 15.475 310.925 15.805 ;
        RECT 310.595 10.035 310.925 10.365 ;
        RECT 310.595 8.675 310.925 9.005 ;
        RECT 310.595 7.315 310.925 7.645 ;
        RECT 310.595 5.955 310.925 6.285 ;
        RECT 310.595 4.595 310.925 4.925 ;
        RECT 310.595 3.235 310.925 3.565 ;
        RECT 310.595 1.875 310.925 2.205 ;
        RECT 310.595 0.515 310.925 0.845 ;
        RECT 310.6 -8.32 310.92 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 311.955 15.475 312.285 15.805 ;
        RECT 311.955 10.035 312.285 10.365 ;
        RECT 311.955 8.675 312.285 9.005 ;
        RECT 311.955 7.315 312.285 7.645 ;
        RECT 311.955 5.955 312.285 6.285 ;
        RECT 311.955 4.595 312.285 4.925 ;
        RECT 311.955 3.235 312.285 3.565 ;
        RECT 311.955 1.875 312.285 2.205 ;
        RECT 311.955 0.515 312.285 0.845 ;
        RECT 311.96 -8.32 312.28 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.315 15.475 313.645 15.805 ;
        RECT 313.315 10.035 313.645 10.365 ;
        RECT 313.315 8.675 313.645 9.005 ;
        RECT 313.315 7.315 313.645 7.645 ;
        RECT 313.315 5.955 313.645 6.285 ;
        RECT 313.315 4.595 313.645 4.925 ;
        RECT 313.315 3.235 313.645 3.565 ;
        RECT 313.315 1.875 313.645 2.205 ;
        RECT 313.315 0.515 313.645 0.845 ;
        RECT 313.32 -8.32 313.64 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 314.675 15.475 315.005 15.805 ;
        RECT 314.675 10.035 315.005 10.365 ;
        RECT 314.675 8.675 315.005 9.005 ;
        RECT 314.675 7.315 315.005 7.645 ;
        RECT 314.675 5.955 315.005 6.285 ;
        RECT 314.675 4.595 315.005 4.925 ;
        RECT 314.675 3.235 315.005 3.565 ;
        RECT 314.675 1.875 315.005 2.205 ;
        RECT 314.675 0.515 315.005 0.845 ;
        RECT 314.68 -8.32 315 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 316.035 15.475 316.365 15.805 ;
        RECT 316.035 11.395 316.365 11.725 ;
        RECT 316.035 10.035 316.365 10.365 ;
        RECT 316.035 8.675 316.365 9.005 ;
        RECT 316.035 7.315 316.365 7.645 ;
        RECT 316.035 5.955 316.365 6.285 ;
        RECT 316.035 4.595 316.365 4.925 ;
        RECT 316.035 3.235 316.365 3.565 ;
        RECT 316.035 1.875 316.365 2.205 ;
        RECT 316.035 0.515 316.365 0.845 ;
        RECT 316.04 -8.32 316.36 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 317.395 15.475 317.725 15.805 ;
        RECT 317.395 11.395 317.725 11.725 ;
        RECT 317.395 10.035 317.725 10.365 ;
        RECT 317.395 8.675 317.725 9.005 ;
        RECT 317.395 7.315 317.725 7.645 ;
        RECT 317.395 5.955 317.725 6.285 ;
        RECT 317.395 4.595 317.725 4.925 ;
        RECT 317.395 3.235 317.725 3.565 ;
        RECT 317.395 1.875 317.725 2.205 ;
        RECT 317.395 0.515 317.725 0.845 ;
        RECT 317.4 -8.32 317.72 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.755 15.475 319.085 15.805 ;
        RECT 318.755 11.395 319.085 11.725 ;
        RECT 318.755 10.035 319.085 10.365 ;
        RECT 318.755 8.675 319.085 9.005 ;
        RECT 318.755 7.315 319.085 7.645 ;
        RECT 318.755 5.955 319.085 6.285 ;
        RECT 318.755 4.595 319.085 4.925 ;
        RECT 318.755 3.235 319.085 3.565 ;
        RECT 318.755 1.875 319.085 2.205 ;
        RECT 318.755 0.515 319.085 0.845 ;
        RECT 318.76 -8.32 319.08 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 320.115 15.475 320.445 15.805 ;
        RECT 320.115 10.035 320.445 10.365 ;
        RECT 320.115 8.675 320.445 9.005 ;
        RECT 320.115 7.315 320.445 7.645 ;
        RECT 320.115 5.955 320.445 6.285 ;
        RECT 320.115 4.595 320.445 4.925 ;
        RECT 320.115 3.235 320.445 3.565 ;
        RECT 320.115 1.875 320.445 2.205 ;
        RECT 320.115 0.515 320.445 0.845 ;
        RECT 320.12 -8.32 320.44 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 321.475 15.475 321.805 15.805 ;
        RECT 321.475 10.035 321.805 10.365 ;
        RECT 321.475 8.675 321.805 9.005 ;
        RECT 321.475 7.315 321.805 7.645 ;
        RECT 321.475 5.955 321.805 6.285 ;
        RECT 321.475 4.595 321.805 4.925 ;
        RECT 321.475 3.235 321.805 3.565 ;
        RECT 321.475 1.875 321.805 2.205 ;
        RECT 321.475 0.515 321.805 0.845 ;
        RECT 321.48 -8.32 321.8 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 322.835 15.475 323.165 15.805 ;
        RECT 322.835 10.035 323.165 10.365 ;
        RECT 322.835 8.675 323.165 9.005 ;
        RECT 322.835 7.315 323.165 7.645 ;
        RECT 322.835 5.955 323.165 6.285 ;
        RECT 322.835 4.595 323.165 4.925 ;
        RECT 322.835 3.235 323.165 3.565 ;
        RECT 322.835 1.875 323.165 2.205 ;
        RECT 322.835 0.515 323.165 0.845 ;
        RECT 322.84 -8.32 323.16 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.195 15.475 324.525 15.805 ;
        RECT 324.195 10.035 324.525 10.365 ;
        RECT 324.195 8.675 324.525 9.005 ;
        RECT 324.195 7.315 324.525 7.645 ;
        RECT 324.195 5.955 324.525 6.285 ;
        RECT 324.195 4.595 324.525 4.925 ;
        RECT 324.195 3.235 324.525 3.565 ;
        RECT 324.195 1.875 324.525 2.205 ;
        RECT 324.195 0.515 324.525 0.845 ;
        RECT 324.2 -8.32 324.52 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 325.555 15.475 325.885 15.805 ;
        RECT 325.555 10.035 325.885 10.365 ;
        RECT 325.555 8.675 325.885 9.005 ;
        RECT 325.555 7.315 325.885 7.645 ;
        RECT 325.555 5.955 325.885 6.285 ;
        RECT 325.555 4.595 325.885 4.925 ;
        RECT 325.555 3.235 325.885 3.565 ;
        RECT 325.555 1.875 325.885 2.205 ;
        RECT 325.555 0.515 325.885 0.845 ;
        RECT 325.56 -8.32 325.88 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 326.915 15.475 327.245 15.805 ;
        RECT 326.915 11.395 327.245 11.725 ;
        RECT 326.915 10.035 327.245 10.365 ;
        RECT 326.915 8.675 327.245 9.005 ;
        RECT 326.915 7.315 327.245 7.645 ;
        RECT 326.915 5.955 327.245 6.285 ;
        RECT 326.915 4.595 327.245 4.925 ;
        RECT 326.915 3.235 327.245 3.565 ;
        RECT 326.915 1.875 327.245 2.205 ;
        RECT 326.915 0.515 327.245 0.845 ;
        RECT 326.92 -8.32 327.24 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 328.275 15.475 328.605 15.805 ;
        RECT 328.275 11.395 328.605 11.725 ;
        RECT 328.275 10.035 328.605 10.365 ;
        RECT 328.275 8.675 328.605 9.005 ;
        RECT 328.275 7.315 328.605 7.645 ;
        RECT 328.275 5.955 328.605 6.285 ;
        RECT 328.275 4.595 328.605 4.925 ;
        RECT 328.275 3.235 328.605 3.565 ;
        RECT 328.275 1.875 328.605 2.205 ;
        RECT 328.275 0.515 328.605 0.845 ;
        RECT 328.28 -8.32 328.6 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 329.635 15.475 329.965 15.805 ;
        RECT 329.635 11.395 329.965 11.725 ;
        RECT 329.635 10.035 329.965 10.365 ;
        RECT 329.635 8.675 329.965 9.005 ;
        RECT 329.635 7.315 329.965 7.645 ;
        RECT 329.635 5.955 329.965 6.285 ;
        RECT 329.635 4.595 329.965 4.925 ;
        RECT 329.635 3.235 329.965 3.565 ;
        RECT 329.635 1.875 329.965 2.205 ;
        RECT 329.635 0.515 329.965 0.845 ;
        RECT 329.64 -8.32 329.96 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.995 15.475 331.325 15.805 ;
        RECT 330.995 10.035 331.325 10.365 ;
        RECT 330.995 8.675 331.325 9.005 ;
        RECT 330.995 7.315 331.325 7.645 ;
        RECT 330.995 5.955 331.325 6.285 ;
        RECT 330.995 4.595 331.325 4.925 ;
        RECT 330.995 3.235 331.325 3.565 ;
        RECT 330.995 1.875 331.325 2.205 ;
        RECT 330.995 0.515 331.325 0.845 ;
        RECT 331 -8.32 331.32 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 332.355 15.475 332.685 15.805 ;
        RECT 332.355 10.035 332.685 10.365 ;
        RECT 332.355 8.675 332.685 9.005 ;
        RECT 332.355 7.315 332.685 7.645 ;
        RECT 332.355 5.955 332.685 6.285 ;
        RECT 332.355 4.595 332.685 4.925 ;
        RECT 332.355 3.235 332.685 3.565 ;
        RECT 332.355 1.875 332.685 2.205 ;
        RECT 332.355 0.515 332.685 0.845 ;
        RECT 332.36 -8.32 332.68 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 333.715 15.475 334.045 15.805 ;
        RECT 333.715 10.035 334.045 10.365 ;
        RECT 333.715 8.675 334.045 9.005 ;
        RECT 333.715 7.315 334.045 7.645 ;
        RECT 333.715 5.955 334.045 6.285 ;
        RECT 333.715 4.595 334.045 4.925 ;
        RECT 333.715 3.235 334.045 3.565 ;
        RECT 333.715 1.875 334.045 2.205 ;
        RECT 333.715 0.515 334.045 0.845 ;
        RECT 333.72 -8.32 334.04 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.075 15.475 335.405 15.805 ;
        RECT 335.075 10.035 335.405 10.365 ;
        RECT 335.075 8.675 335.405 9.005 ;
        RECT 335.075 7.315 335.405 7.645 ;
        RECT 335.075 5.955 335.405 6.285 ;
        RECT 335.075 4.595 335.405 4.925 ;
        RECT 335.075 3.235 335.405 3.565 ;
        RECT 335.075 1.875 335.405 2.205 ;
        RECT 335.075 0.515 335.405 0.845 ;
        RECT 335.08 -8.32 335.4 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 336.435 15.475 336.765 15.805 ;
        RECT 336.435 10.035 336.765 10.365 ;
        RECT 336.435 8.675 336.765 9.005 ;
        RECT 336.435 7.315 336.765 7.645 ;
        RECT 336.435 5.955 336.765 6.285 ;
        RECT 336.435 4.595 336.765 4.925 ;
        RECT 336.435 3.235 336.765 3.565 ;
        RECT 336.435 1.875 336.765 2.205 ;
        RECT 336.435 0.515 336.765 0.845 ;
        RECT 336.44 -8.32 336.76 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 337.795 15.475 338.125 15.805 ;
        RECT 337.795 10.035 338.125 10.365 ;
        RECT 337.795 8.675 338.125 9.005 ;
        RECT 337.795 7.315 338.125 7.645 ;
        RECT 337.795 5.955 338.125 6.285 ;
        RECT 337.795 4.595 338.125 4.925 ;
        RECT 337.795 3.235 338.125 3.565 ;
        RECT 337.795 1.875 338.125 2.205 ;
        RECT 337.795 0.515 338.125 0.845 ;
        RECT 337.8 -8.32 338.12 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 339.155 15.475 339.485 15.805 ;
        RECT 339.155 11.395 339.485 11.725 ;
        RECT 339.155 10.035 339.485 10.365 ;
        RECT 339.155 8.675 339.485 9.005 ;
        RECT 339.155 7.315 339.485 7.645 ;
        RECT 339.155 5.955 339.485 6.285 ;
        RECT 339.155 4.595 339.485 4.925 ;
        RECT 339.155 3.235 339.485 3.565 ;
        RECT 339.155 1.875 339.485 2.205 ;
        RECT 339.155 0.515 339.485 0.845 ;
        RECT 339.16 -8.32 339.48 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 340.515 15.475 340.845 15.805 ;
        RECT 340.515 11.395 340.845 11.725 ;
        RECT 340.515 10.035 340.845 10.365 ;
        RECT 340.515 8.675 340.845 9.005 ;
        RECT 340.515 7.315 340.845 7.645 ;
        RECT 340.515 5.955 340.845 6.285 ;
        RECT 340.515 4.595 340.845 4.925 ;
        RECT 340.515 3.235 340.845 3.565 ;
        RECT 340.515 1.875 340.845 2.205 ;
        RECT 340.515 0.515 340.845 0.845 ;
        RECT 340.52 -8.32 340.84 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 341.875 15.475 342.205 15.805 ;
        RECT 341.875 11.395 342.205 11.725 ;
        RECT 341.875 10.035 342.205 10.365 ;
        RECT 341.875 8.675 342.205 9.005 ;
        RECT 341.875 7.315 342.205 7.645 ;
        RECT 341.875 5.955 342.205 6.285 ;
        RECT 341.875 4.595 342.205 4.925 ;
        RECT 341.875 3.235 342.205 3.565 ;
        RECT 341.875 1.875 342.205 2.205 ;
        RECT 341.875 0.515 342.205 0.845 ;
        RECT 341.88 -8.32 342.2 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 343.235 15.475 343.565 15.805 ;
        RECT 343.235 10.035 343.565 10.365 ;
        RECT 343.235 8.675 343.565 9.005 ;
        RECT 343.235 7.315 343.565 7.645 ;
        RECT 343.235 5.955 343.565 6.285 ;
        RECT 343.235 4.595 343.565 4.925 ;
        RECT 343.235 3.235 343.565 3.565 ;
        RECT 343.235 1.875 343.565 2.205 ;
        RECT 343.235 0.515 343.565 0.845 ;
        RECT 343.24 -8.32 343.56 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 344.595 15.475 344.925 15.805 ;
        RECT 344.595 10.035 344.925 10.365 ;
        RECT 344.595 8.675 344.925 9.005 ;
        RECT 344.595 7.315 344.925 7.645 ;
        RECT 344.595 5.955 344.925 6.285 ;
        RECT 344.595 4.595 344.925 4.925 ;
        RECT 344.595 3.235 344.925 3.565 ;
        RECT 344.595 1.875 344.925 2.205 ;
        RECT 344.595 0.515 344.925 0.845 ;
        RECT 344.6 -8.32 344.92 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 345.955 15.475 346.285 15.805 ;
        RECT 345.955 10.035 346.285 10.365 ;
        RECT 345.955 8.675 346.285 9.005 ;
        RECT 345.955 7.315 346.285 7.645 ;
        RECT 345.955 5.955 346.285 6.285 ;
        RECT 345.955 4.595 346.285 4.925 ;
        RECT 345.955 3.235 346.285 3.565 ;
        RECT 345.955 1.875 346.285 2.205 ;
        RECT 345.955 0.515 346.285 0.845 ;
        RECT 345.96 -8.32 346.28 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 347.315 15.475 347.645 15.805 ;
        RECT 347.315 10.035 347.645 10.365 ;
        RECT 347.315 8.675 347.645 9.005 ;
        RECT 347.315 7.315 347.645 7.645 ;
        RECT 347.315 5.955 347.645 6.285 ;
        RECT 347.315 4.595 347.645 4.925 ;
        RECT 347.315 3.235 347.645 3.565 ;
        RECT 347.315 1.875 347.645 2.205 ;
        RECT 347.315 0.515 347.645 0.845 ;
        RECT 347.32 -8.32 347.64 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 348.675 15.475 349.005 15.805 ;
        RECT 348.675 10.035 349.005 10.365 ;
        RECT 348.675 8.675 349.005 9.005 ;
        RECT 348.675 7.315 349.005 7.645 ;
        RECT 348.675 5.955 349.005 6.285 ;
        RECT 348.675 4.595 349.005 4.925 ;
        RECT 348.675 3.235 349.005 3.565 ;
        RECT 348.675 1.875 349.005 2.205 ;
        RECT 348.675 0.515 349.005 0.845 ;
        RECT 348.68 -8.32 349 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 350.035 15.475 350.365 15.805 ;
        RECT 350.035 10.035 350.365 10.365 ;
        RECT 350.035 8.675 350.365 9.005 ;
        RECT 350.035 7.315 350.365 7.645 ;
        RECT 350.035 5.955 350.365 6.285 ;
        RECT 350.035 4.595 350.365 4.925 ;
        RECT 350.035 3.235 350.365 3.565 ;
        RECT 350.035 1.875 350.365 2.205 ;
        RECT 350.035 0.515 350.365 0.845 ;
        RECT 350.04 -8.32 350.36 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 351.395 15.475 351.725 15.805 ;
        RECT 351.395 11.395 351.725 11.725 ;
        RECT 351.395 10.035 351.725 10.365 ;
        RECT 351.395 8.675 351.725 9.005 ;
        RECT 351.395 7.315 351.725 7.645 ;
        RECT 351.395 5.955 351.725 6.285 ;
        RECT 351.395 4.595 351.725 4.925 ;
        RECT 351.395 3.235 351.725 3.565 ;
        RECT 351.395 1.875 351.725 2.205 ;
        RECT 351.395 0.515 351.725 0.845 ;
        RECT 351.4 -8.32 351.72 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 352.755 15.475 353.085 15.805 ;
        RECT 352.755 11.395 353.085 11.725 ;
        RECT 352.755 10.035 353.085 10.365 ;
        RECT 352.755 8.675 353.085 9.005 ;
        RECT 352.755 7.315 353.085 7.645 ;
        RECT 352.755 5.955 353.085 6.285 ;
        RECT 352.755 4.595 353.085 4.925 ;
        RECT 352.755 3.235 353.085 3.565 ;
        RECT 352.755 1.875 353.085 2.205 ;
        RECT 352.755 0.515 353.085 0.845 ;
        RECT 352.76 -8.32 353.08 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.115 15.475 354.445 15.805 ;
        RECT 354.115 11.395 354.445 11.725 ;
        RECT 354.115 10.035 354.445 10.365 ;
        RECT 354.115 8.675 354.445 9.005 ;
        RECT 354.115 7.315 354.445 7.645 ;
        RECT 354.115 5.955 354.445 6.285 ;
        RECT 354.115 4.595 354.445 4.925 ;
        RECT 354.115 3.235 354.445 3.565 ;
        RECT 354.115 1.875 354.445 2.205 ;
        RECT 354.115 0.515 354.445 0.845 ;
        RECT 354.12 -8.32 354.44 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 355.475 15.475 355.805 15.805 ;
        RECT 355.475 10.035 355.805 10.365 ;
        RECT 355.475 8.675 355.805 9.005 ;
        RECT 355.475 7.315 355.805 7.645 ;
        RECT 355.475 5.955 355.805 6.285 ;
        RECT 355.475 4.595 355.805 4.925 ;
        RECT 355.475 3.235 355.805 3.565 ;
        RECT 355.475 1.875 355.805 2.205 ;
        RECT 355.475 0.515 355.805 0.845 ;
        RECT 355.48 -8.32 355.8 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 356.835 15.475 357.165 15.805 ;
        RECT 356.835 10.035 357.165 10.365 ;
        RECT 356.835 8.675 357.165 9.005 ;
        RECT 356.835 7.315 357.165 7.645 ;
        RECT 356.835 5.955 357.165 6.285 ;
        RECT 356.835 4.595 357.165 4.925 ;
        RECT 356.835 3.235 357.165 3.565 ;
        RECT 356.835 1.875 357.165 2.205 ;
        RECT 356.835 0.515 357.165 0.845 ;
        RECT 356.84 -8.32 357.16 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 358.195 15.475 358.525 15.805 ;
        RECT 358.195 10.035 358.525 10.365 ;
        RECT 358.195 8.675 358.525 9.005 ;
        RECT 358.195 7.315 358.525 7.645 ;
        RECT 358.195 5.955 358.525 6.285 ;
        RECT 358.195 4.595 358.525 4.925 ;
        RECT 358.195 3.235 358.525 3.565 ;
        RECT 358.195 1.875 358.525 2.205 ;
        RECT 358.195 0.515 358.525 0.845 ;
        RECT 358.2 -8.32 358.52 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 359.555 15.475 359.885 15.805 ;
        RECT 359.555 10.035 359.885 10.365 ;
        RECT 359.555 8.675 359.885 9.005 ;
        RECT 359.555 7.315 359.885 7.645 ;
        RECT 359.555 5.955 359.885 6.285 ;
        RECT 359.555 4.595 359.885 4.925 ;
        RECT 359.555 3.235 359.885 3.565 ;
        RECT 359.555 1.875 359.885 2.205 ;
        RECT 359.555 0.515 359.885 0.845 ;
        RECT 359.56 -8.32 359.88 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 360.915 15.475 361.245 15.805 ;
        RECT 360.915 10.035 361.245 10.365 ;
        RECT 360.915 8.675 361.245 9.005 ;
        RECT 360.915 7.315 361.245 7.645 ;
        RECT 360.915 5.955 361.245 6.285 ;
        RECT 360.915 4.595 361.245 4.925 ;
        RECT 360.915 3.235 361.245 3.565 ;
        RECT 360.915 1.875 361.245 2.205 ;
        RECT 360.915 0.515 361.245 0.845 ;
        RECT 360.92 -8.32 361.24 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 362.275 15.475 362.605 15.805 ;
        RECT 362.275 10.035 362.605 10.365 ;
        RECT 362.275 8.675 362.605 9.005 ;
        RECT 362.275 7.315 362.605 7.645 ;
        RECT 362.275 5.955 362.605 6.285 ;
        RECT 362.275 4.595 362.605 4.925 ;
        RECT 362.275 3.235 362.605 3.565 ;
        RECT 362.275 1.875 362.605 2.205 ;
        RECT 362.275 0.515 362.605 0.845 ;
        RECT 362.28 -8.32 362.6 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 363.635 15.475 363.965 15.805 ;
        RECT 363.635 11.395 363.965 11.725 ;
        RECT 363.635 10.035 363.965 10.365 ;
        RECT 363.635 8.675 363.965 9.005 ;
        RECT 363.635 7.315 363.965 7.645 ;
        RECT 363.635 5.955 363.965 6.285 ;
        RECT 363.635 4.595 363.965 4.925 ;
        RECT 363.635 3.235 363.965 3.565 ;
        RECT 363.635 1.875 363.965 2.205 ;
        RECT 363.635 0.515 363.965 0.845 ;
        RECT 363.64 -8.32 363.96 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 364.995 15.475 365.325 15.805 ;
        RECT 364.995 11.395 365.325 11.725 ;
        RECT 364.995 10.035 365.325 10.365 ;
        RECT 364.995 8.675 365.325 9.005 ;
        RECT 364.995 7.315 365.325 7.645 ;
        RECT 364.995 5.955 365.325 6.285 ;
        RECT 364.995 4.595 365.325 4.925 ;
        RECT 364.995 3.235 365.325 3.565 ;
        RECT 364.995 1.875 365.325 2.205 ;
        RECT 364.995 0.515 365.325 0.845 ;
        RECT 365 -8.32 365.32 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 366.355 15.475 366.685 15.805 ;
        RECT 366.355 11.395 366.685 11.725 ;
        RECT 366.355 10.035 366.685 10.365 ;
        RECT 366.355 8.675 366.685 9.005 ;
        RECT 366.355 7.315 366.685 7.645 ;
        RECT 366.355 5.955 366.685 6.285 ;
        RECT 366.355 4.595 366.685 4.925 ;
        RECT 366.355 3.235 366.685 3.565 ;
        RECT 366.355 1.875 366.685 2.205 ;
        RECT 366.355 0.515 366.685 0.845 ;
        RECT 366.36 -8.32 366.68 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 367.715 15.475 368.045 15.805 ;
        RECT 367.715 10.035 368.045 10.365 ;
        RECT 367.715 8.675 368.045 9.005 ;
        RECT 367.715 7.315 368.045 7.645 ;
        RECT 367.715 5.955 368.045 6.285 ;
        RECT 367.715 4.595 368.045 4.925 ;
        RECT 367.715 3.235 368.045 3.565 ;
        RECT 367.715 1.875 368.045 2.205 ;
        RECT 367.715 0.515 368.045 0.845 ;
        RECT 367.72 -8.32 368.04 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 369.075 15.475 369.405 15.805 ;
        RECT 369.075 10.035 369.405 10.365 ;
        RECT 369.075 8.675 369.405 9.005 ;
        RECT 369.075 7.315 369.405 7.645 ;
        RECT 369.075 5.955 369.405 6.285 ;
        RECT 369.075 4.595 369.405 4.925 ;
        RECT 369.075 3.235 369.405 3.565 ;
        RECT 369.075 1.875 369.405 2.205 ;
        RECT 369.075 0.515 369.405 0.845 ;
        RECT 369.08 -8.32 369.4 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 370.435 15.475 370.765 15.805 ;
        RECT 370.435 10.035 370.765 10.365 ;
        RECT 370.435 8.675 370.765 9.005 ;
        RECT 370.435 7.315 370.765 7.645 ;
        RECT 370.435 5.955 370.765 6.285 ;
        RECT 370.435 4.595 370.765 4.925 ;
        RECT 370.435 3.235 370.765 3.565 ;
        RECT 370.435 1.875 370.765 2.205 ;
        RECT 370.435 0.515 370.765 0.845 ;
        RECT 370.44 -8.32 370.76 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 371.795 15.475 372.125 15.805 ;
        RECT 371.795 10.035 372.125 10.365 ;
        RECT 371.795 8.675 372.125 9.005 ;
        RECT 371.795 7.315 372.125 7.645 ;
        RECT 371.795 5.955 372.125 6.285 ;
        RECT 371.795 4.595 372.125 4.925 ;
        RECT 371.795 3.235 372.125 3.565 ;
        RECT 371.795 1.875 372.125 2.205 ;
        RECT 371.795 0.515 372.125 0.845 ;
        RECT 371.8 -8.32 372.12 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 373.155 15.475 373.485 15.805 ;
        RECT 373.155 10.035 373.485 10.365 ;
        RECT 373.155 8.675 373.485 9.005 ;
        RECT 373.155 7.315 373.485 7.645 ;
        RECT 373.155 5.955 373.485 6.285 ;
        RECT 373.155 4.595 373.485 4.925 ;
        RECT 373.155 3.235 373.485 3.565 ;
        RECT 373.155 1.875 373.485 2.205 ;
        RECT 373.155 0.515 373.485 0.845 ;
        RECT 373.16 -8.32 373.48 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 374.515 15.475 374.845 15.805 ;
        RECT 374.515 10.035 374.845 10.365 ;
        RECT 374.515 8.675 374.845 9.005 ;
        RECT 374.515 7.315 374.845 7.645 ;
        RECT 374.515 5.955 374.845 6.285 ;
        RECT 374.515 4.595 374.845 4.925 ;
        RECT 374.515 3.235 374.845 3.565 ;
        RECT 374.515 1.875 374.845 2.205 ;
        RECT 374.515 0.515 374.845 0.845 ;
        RECT 374.52 -8.32 374.84 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 375.875 11.395 376.205 11.725 ;
        RECT 375.875 10.035 376.205 10.365 ;
        RECT 375.875 8.675 376.205 9.005 ;
        RECT 375.875 7.315 376.205 7.645 ;
        RECT 375.875 5.955 376.205 6.285 ;
        RECT 375.875 4.595 376.205 4.925 ;
        RECT 375.875 3.235 376.205 3.565 ;
        RECT 375.875 1.875 376.205 2.205 ;
        RECT 375.875 0.515 376.205 0.845 ;
        RECT 375.88 -8.32 376.2 15.805 ;
        RECT 375.875 15.475 376.205 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.755 15.475 115.085 15.805 ;
        RECT 114.755 11.395 115.085 11.725 ;
        RECT 114.755 10.035 115.085 10.365 ;
        RECT 114.755 8.675 115.085 9.005 ;
        RECT 114.755 7.315 115.085 7.645 ;
        RECT 114.755 5.955 115.085 6.285 ;
        RECT 114.755 4.595 115.085 4.925 ;
        RECT 114.755 3.235 115.085 3.565 ;
        RECT 114.755 1.875 115.085 2.205 ;
        RECT 114.755 0.515 115.085 0.845 ;
        RECT 114.76 -8.32 115.08 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.115 15.475 116.445 15.805 ;
        RECT 116.115 10.035 116.445 10.365 ;
        RECT 116.115 8.675 116.445 9.005 ;
        RECT 116.115 7.315 116.445 7.645 ;
        RECT 116.115 5.955 116.445 6.285 ;
        RECT 116.115 4.595 116.445 4.925 ;
        RECT 116.115 3.235 116.445 3.565 ;
        RECT 116.115 1.875 116.445 2.205 ;
        RECT 116.115 0.515 116.445 0.845 ;
        RECT 116.12 -8.32 116.44 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 117.475 15.475 117.805 15.805 ;
        RECT 117.475 10.035 117.805 10.365 ;
        RECT 117.475 8.675 117.805 9.005 ;
        RECT 117.475 7.315 117.805 7.645 ;
        RECT 117.475 5.955 117.805 6.285 ;
        RECT 117.475 4.595 117.805 4.925 ;
        RECT 117.475 3.235 117.805 3.565 ;
        RECT 117.475 1.875 117.805 2.205 ;
        RECT 117.475 0.515 117.805 0.845 ;
        RECT 117.48 -8.32 117.8 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.835 15.475 119.165 15.805 ;
        RECT 118.835 10.035 119.165 10.365 ;
        RECT 118.835 8.675 119.165 9.005 ;
        RECT 118.835 7.315 119.165 7.645 ;
        RECT 118.835 5.955 119.165 6.285 ;
        RECT 118.835 4.595 119.165 4.925 ;
        RECT 118.835 3.235 119.165 3.565 ;
        RECT 118.835 1.875 119.165 2.205 ;
        RECT 118.835 0.515 119.165 0.845 ;
        RECT 118.84 -8.32 119.16 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.195 15.475 120.525 15.805 ;
        RECT 120.195 10.035 120.525 10.365 ;
        RECT 120.195 8.675 120.525 9.005 ;
        RECT 120.195 7.315 120.525 7.645 ;
        RECT 120.195 5.955 120.525 6.285 ;
        RECT 120.195 4.595 120.525 4.925 ;
        RECT 120.195 3.235 120.525 3.565 ;
        RECT 120.195 1.875 120.525 2.205 ;
        RECT 120.195 0.515 120.525 0.845 ;
        RECT 120.2 -8.32 120.52 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 121.555 15.475 121.885 15.805 ;
        RECT 121.555 10.035 121.885 10.365 ;
        RECT 121.555 8.675 121.885 9.005 ;
        RECT 121.555 7.315 121.885 7.645 ;
        RECT 121.555 5.955 121.885 6.285 ;
        RECT 121.555 4.595 121.885 4.925 ;
        RECT 121.555 3.235 121.885 3.565 ;
        RECT 121.555 1.875 121.885 2.205 ;
        RECT 121.555 0.515 121.885 0.845 ;
        RECT 121.56 -8.32 121.88 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.915 15.475 123.245 15.805 ;
        RECT 122.915 11.395 123.245 11.725 ;
        RECT 122.915 10.035 123.245 10.365 ;
        RECT 122.915 8.675 123.245 9.005 ;
        RECT 122.915 7.315 123.245 7.645 ;
        RECT 122.915 5.955 123.245 6.285 ;
        RECT 122.915 4.595 123.245 4.925 ;
        RECT 122.915 3.235 123.245 3.565 ;
        RECT 122.915 1.875 123.245 2.205 ;
        RECT 122.915 0.515 123.245 0.845 ;
        RECT 122.92 -8.32 123.24 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.275 15.475 124.605 15.805 ;
        RECT 124.275 11.395 124.605 11.725 ;
        RECT 124.275 10.035 124.605 10.365 ;
        RECT 124.275 8.675 124.605 9.005 ;
        RECT 124.275 7.315 124.605 7.645 ;
        RECT 124.275 5.955 124.605 6.285 ;
        RECT 124.275 4.595 124.605 4.925 ;
        RECT 124.275 3.235 124.605 3.565 ;
        RECT 124.275 1.875 124.605 2.205 ;
        RECT 124.275 0.515 124.605 0.845 ;
        RECT 124.28 -8.32 124.6 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.635 15.475 125.965 15.805 ;
        RECT 125.635 11.395 125.965 11.725 ;
        RECT 125.635 10.035 125.965 10.365 ;
        RECT 125.635 8.675 125.965 9.005 ;
        RECT 125.635 7.315 125.965 7.645 ;
        RECT 125.635 5.955 125.965 6.285 ;
        RECT 125.635 4.595 125.965 4.925 ;
        RECT 125.635 3.235 125.965 3.565 ;
        RECT 125.635 1.875 125.965 2.205 ;
        RECT 125.635 0.515 125.965 0.845 ;
        RECT 125.64 -8.32 125.96 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.995 15.475 127.325 15.805 ;
        RECT 126.995 10.035 127.325 10.365 ;
        RECT 126.995 8.675 127.325 9.005 ;
        RECT 126.995 7.315 127.325 7.645 ;
        RECT 126.995 5.955 127.325 6.285 ;
        RECT 126.995 4.595 127.325 4.925 ;
        RECT 126.995 3.235 127.325 3.565 ;
        RECT 126.995 1.875 127.325 2.205 ;
        RECT 126.995 0.515 127.325 0.845 ;
        RECT 127 -8.32 127.32 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.355 15.475 128.685 15.805 ;
        RECT 128.355 10.035 128.685 10.365 ;
        RECT 128.355 8.675 128.685 9.005 ;
        RECT 128.355 7.315 128.685 7.645 ;
        RECT 128.355 5.955 128.685 6.285 ;
        RECT 128.355 4.595 128.685 4.925 ;
        RECT 128.355 3.235 128.685 3.565 ;
        RECT 128.355 1.875 128.685 2.205 ;
        RECT 128.355 0.515 128.685 0.845 ;
        RECT 128.36 -8.32 128.68 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.715 15.475 130.045 15.805 ;
        RECT 129.715 10.035 130.045 10.365 ;
        RECT 129.715 8.675 130.045 9.005 ;
        RECT 129.715 7.315 130.045 7.645 ;
        RECT 129.715 5.955 130.045 6.285 ;
        RECT 129.715 4.595 130.045 4.925 ;
        RECT 129.715 3.235 130.045 3.565 ;
        RECT 129.715 1.875 130.045 2.205 ;
        RECT 129.715 0.515 130.045 0.845 ;
        RECT 129.72 -8.32 130.04 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.075 15.475 131.405 15.805 ;
        RECT 131.075 10.035 131.405 10.365 ;
        RECT 131.075 8.675 131.405 9.005 ;
        RECT 131.075 7.315 131.405 7.645 ;
        RECT 131.075 5.955 131.405 6.285 ;
        RECT 131.075 4.595 131.405 4.925 ;
        RECT 131.075 3.235 131.405 3.565 ;
        RECT 131.075 1.875 131.405 2.205 ;
        RECT 131.075 0.515 131.405 0.845 ;
        RECT 131.08 -8.32 131.4 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.435 15.475 132.765 15.805 ;
        RECT 132.435 10.035 132.765 10.365 ;
        RECT 132.435 8.675 132.765 9.005 ;
        RECT 132.435 7.315 132.765 7.645 ;
        RECT 132.435 5.955 132.765 6.285 ;
        RECT 132.435 4.595 132.765 4.925 ;
        RECT 132.435 3.235 132.765 3.565 ;
        RECT 132.435 1.875 132.765 2.205 ;
        RECT 132.435 0.515 132.765 0.845 ;
        RECT 132.44 -8.32 132.76 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.795 15.475 134.125 15.805 ;
        RECT 133.795 10.035 134.125 10.365 ;
        RECT 133.795 8.675 134.125 9.005 ;
        RECT 133.795 7.315 134.125 7.645 ;
        RECT 133.795 5.955 134.125 6.285 ;
        RECT 133.795 4.595 134.125 4.925 ;
        RECT 133.795 3.235 134.125 3.565 ;
        RECT 133.795 1.875 134.125 2.205 ;
        RECT 133.795 0.515 134.125 0.845 ;
        RECT 133.8 -8.32 134.12 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.155 15.475 135.485 15.805 ;
        RECT 135.155 11.395 135.485 11.725 ;
        RECT 135.155 10.035 135.485 10.365 ;
        RECT 135.155 8.675 135.485 9.005 ;
        RECT 135.155 7.315 135.485 7.645 ;
        RECT 135.155 5.955 135.485 6.285 ;
        RECT 135.155 4.595 135.485 4.925 ;
        RECT 135.155 3.235 135.485 3.565 ;
        RECT 135.155 1.875 135.485 2.205 ;
        RECT 135.155 0.515 135.485 0.845 ;
        RECT 135.16 -8.32 135.48 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 136.515 15.475 136.845 15.805 ;
        RECT 136.515 11.395 136.845 11.725 ;
        RECT 136.515 10.035 136.845 10.365 ;
        RECT 136.515 8.675 136.845 9.005 ;
        RECT 136.515 7.315 136.845 7.645 ;
        RECT 136.515 5.955 136.845 6.285 ;
        RECT 136.515 4.595 136.845 4.925 ;
        RECT 136.515 3.235 136.845 3.565 ;
        RECT 136.515 1.875 136.845 2.205 ;
        RECT 136.515 0.515 136.845 0.845 ;
        RECT 136.52 -8.32 136.84 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.875 15.475 138.205 15.805 ;
        RECT 137.875 11.395 138.205 11.725 ;
        RECT 137.875 10.035 138.205 10.365 ;
        RECT 137.875 8.675 138.205 9.005 ;
        RECT 137.875 7.315 138.205 7.645 ;
        RECT 137.875 5.955 138.205 6.285 ;
        RECT 137.875 4.595 138.205 4.925 ;
        RECT 137.875 3.235 138.205 3.565 ;
        RECT 137.875 1.875 138.205 2.205 ;
        RECT 137.875 0.515 138.205 0.845 ;
        RECT 137.88 -8.32 138.2 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.235 15.475 139.565 15.805 ;
        RECT 139.235 10.035 139.565 10.365 ;
        RECT 139.235 8.675 139.565 9.005 ;
        RECT 139.235 7.315 139.565 7.645 ;
        RECT 139.235 5.955 139.565 6.285 ;
        RECT 139.235 4.595 139.565 4.925 ;
        RECT 139.235 3.235 139.565 3.565 ;
        RECT 139.235 1.875 139.565 2.205 ;
        RECT 139.235 0.515 139.565 0.845 ;
        RECT 139.24 -8.32 139.56 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.595 15.475 140.925 15.805 ;
        RECT 140.595 10.035 140.925 10.365 ;
        RECT 140.595 8.675 140.925 9.005 ;
        RECT 140.595 7.315 140.925 7.645 ;
        RECT 140.595 5.955 140.925 6.285 ;
        RECT 140.595 4.595 140.925 4.925 ;
        RECT 140.595 3.235 140.925 3.565 ;
        RECT 140.595 1.875 140.925 2.205 ;
        RECT 140.595 0.515 140.925 0.845 ;
        RECT 140.6 -8.32 140.92 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.955 15.475 142.285 15.805 ;
        RECT 141.955 10.035 142.285 10.365 ;
        RECT 141.955 8.675 142.285 9.005 ;
        RECT 141.955 7.315 142.285 7.645 ;
        RECT 141.955 5.955 142.285 6.285 ;
        RECT 141.955 4.595 142.285 4.925 ;
        RECT 141.955 3.235 142.285 3.565 ;
        RECT 141.955 1.875 142.285 2.205 ;
        RECT 141.955 0.515 142.285 0.845 ;
        RECT 141.96 -8.32 142.28 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.315 15.475 143.645 15.805 ;
        RECT 143.315 10.035 143.645 10.365 ;
        RECT 143.315 8.675 143.645 9.005 ;
        RECT 143.315 7.315 143.645 7.645 ;
        RECT 143.315 5.955 143.645 6.285 ;
        RECT 143.315 4.595 143.645 4.925 ;
        RECT 143.315 3.235 143.645 3.565 ;
        RECT 143.315 1.875 143.645 2.205 ;
        RECT 143.315 0.515 143.645 0.845 ;
        RECT 143.32 -8.32 143.64 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 144.675 15.475 145.005 15.805 ;
        RECT 144.675 10.035 145.005 10.365 ;
        RECT 144.675 8.675 145.005 9.005 ;
        RECT 144.675 7.315 145.005 7.645 ;
        RECT 144.675 5.955 145.005 6.285 ;
        RECT 144.675 4.595 145.005 4.925 ;
        RECT 144.675 3.235 145.005 3.565 ;
        RECT 144.675 1.875 145.005 2.205 ;
        RECT 144.675 0.515 145.005 0.845 ;
        RECT 144.68 -8.32 145 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.035 15.475 146.365 15.805 ;
        RECT 146.035 10.035 146.365 10.365 ;
        RECT 146.035 8.675 146.365 9.005 ;
        RECT 146.035 7.315 146.365 7.645 ;
        RECT 146.035 5.955 146.365 6.285 ;
        RECT 146.035 4.595 146.365 4.925 ;
        RECT 146.035 3.235 146.365 3.565 ;
        RECT 146.035 1.875 146.365 2.205 ;
        RECT 146.035 0.515 146.365 0.845 ;
        RECT 146.04 -8.32 146.36 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.395 15.475 147.725 15.805 ;
        RECT 147.395 11.395 147.725 11.725 ;
        RECT 147.395 10.035 147.725 10.365 ;
        RECT 147.395 8.675 147.725 9.005 ;
        RECT 147.395 7.315 147.725 7.645 ;
        RECT 147.395 5.955 147.725 6.285 ;
        RECT 147.395 4.595 147.725 4.925 ;
        RECT 147.395 3.235 147.725 3.565 ;
        RECT 147.395 1.875 147.725 2.205 ;
        RECT 147.395 0.515 147.725 0.845 ;
        RECT 147.4 -8.32 147.72 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.755 15.475 149.085 15.805 ;
        RECT 148.755 11.395 149.085 11.725 ;
        RECT 148.755 10.035 149.085 10.365 ;
        RECT 148.755 8.675 149.085 9.005 ;
        RECT 148.755 7.315 149.085 7.645 ;
        RECT 148.755 5.955 149.085 6.285 ;
        RECT 148.755 4.595 149.085 4.925 ;
        RECT 148.755 3.235 149.085 3.565 ;
        RECT 148.755 1.875 149.085 2.205 ;
        RECT 148.755 0.515 149.085 0.845 ;
        RECT 148.76 -8.32 149.08 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.115 15.475 150.445 15.805 ;
        RECT 150.115 11.395 150.445 11.725 ;
        RECT 150.115 10.035 150.445 10.365 ;
        RECT 150.115 8.675 150.445 9.005 ;
        RECT 150.115 7.315 150.445 7.645 ;
        RECT 150.115 5.955 150.445 6.285 ;
        RECT 150.115 4.595 150.445 4.925 ;
        RECT 150.115 3.235 150.445 3.565 ;
        RECT 150.115 1.875 150.445 2.205 ;
        RECT 150.115 0.515 150.445 0.845 ;
        RECT 150.12 -8.32 150.44 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 151.475 15.475 151.805 15.805 ;
        RECT 151.475 10.035 151.805 10.365 ;
        RECT 151.475 8.675 151.805 9.005 ;
        RECT 151.475 7.315 151.805 7.645 ;
        RECT 151.475 5.955 151.805 6.285 ;
        RECT 151.475 4.595 151.805 4.925 ;
        RECT 151.475 3.235 151.805 3.565 ;
        RECT 151.475 1.875 151.805 2.205 ;
        RECT 151.475 0.515 151.805 0.845 ;
        RECT 151.48 -8.32 151.8 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.835 15.475 153.165 15.805 ;
        RECT 152.835 10.035 153.165 10.365 ;
        RECT 152.835 8.675 153.165 9.005 ;
        RECT 152.835 7.315 153.165 7.645 ;
        RECT 152.835 5.955 153.165 6.285 ;
        RECT 152.835 4.595 153.165 4.925 ;
        RECT 152.835 3.235 153.165 3.565 ;
        RECT 152.835 1.875 153.165 2.205 ;
        RECT 152.835 0.515 153.165 0.845 ;
        RECT 152.84 -8.32 153.16 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.195 15.475 154.525 15.805 ;
        RECT 154.195 10.035 154.525 10.365 ;
        RECT 154.195 8.675 154.525 9.005 ;
        RECT 154.195 7.315 154.525 7.645 ;
        RECT 154.195 5.955 154.525 6.285 ;
        RECT 154.195 4.595 154.525 4.925 ;
        RECT 154.195 3.235 154.525 3.565 ;
        RECT 154.195 1.875 154.525 2.205 ;
        RECT 154.195 0.515 154.525 0.845 ;
        RECT 154.2 -8.32 154.52 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.555 15.475 155.885 15.805 ;
        RECT 155.555 10.035 155.885 10.365 ;
        RECT 155.555 8.675 155.885 9.005 ;
        RECT 155.555 7.315 155.885 7.645 ;
        RECT 155.555 5.955 155.885 6.285 ;
        RECT 155.555 4.595 155.885 4.925 ;
        RECT 155.555 3.235 155.885 3.565 ;
        RECT 155.555 1.875 155.885 2.205 ;
        RECT 155.555 0.515 155.885 0.845 ;
        RECT 155.56 -8.32 155.88 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.915 15.475 157.245 15.805 ;
        RECT 156.915 10.035 157.245 10.365 ;
        RECT 156.915 8.675 157.245 9.005 ;
        RECT 156.915 7.315 157.245 7.645 ;
        RECT 156.915 5.955 157.245 6.285 ;
        RECT 156.915 4.595 157.245 4.925 ;
        RECT 156.915 3.235 157.245 3.565 ;
        RECT 156.915 1.875 157.245 2.205 ;
        RECT 156.915 0.515 157.245 0.845 ;
        RECT 156.92 -8.32 157.24 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.275 15.475 158.605 15.805 ;
        RECT 158.275 10.035 158.605 10.365 ;
        RECT 158.275 8.675 158.605 9.005 ;
        RECT 158.275 7.315 158.605 7.645 ;
        RECT 158.275 5.955 158.605 6.285 ;
        RECT 158.275 4.595 158.605 4.925 ;
        RECT 158.275 3.235 158.605 3.565 ;
        RECT 158.275 1.875 158.605 2.205 ;
        RECT 158.275 0.515 158.605 0.845 ;
        RECT 158.28 -8.32 158.6 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.635 15.475 159.965 15.805 ;
        RECT 159.635 11.395 159.965 11.725 ;
        RECT 159.635 10.035 159.965 10.365 ;
        RECT 159.635 8.675 159.965 9.005 ;
        RECT 159.635 7.315 159.965 7.645 ;
        RECT 159.635 5.955 159.965 6.285 ;
        RECT 159.635 4.595 159.965 4.925 ;
        RECT 159.635 3.235 159.965 3.565 ;
        RECT 159.635 1.875 159.965 2.205 ;
        RECT 159.635 0.515 159.965 0.845 ;
        RECT 159.64 -8.32 159.96 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.995 15.475 161.325 15.805 ;
        RECT 160.995 11.395 161.325 11.725 ;
        RECT 160.995 10.035 161.325 10.365 ;
        RECT 160.995 8.675 161.325 9.005 ;
        RECT 160.995 7.315 161.325 7.645 ;
        RECT 160.995 5.955 161.325 6.285 ;
        RECT 160.995 4.595 161.325 4.925 ;
        RECT 160.995 3.235 161.325 3.565 ;
        RECT 160.995 1.875 161.325 2.205 ;
        RECT 160.995 0.515 161.325 0.845 ;
        RECT 161 -8.32 161.32 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 162.355 15.475 162.685 15.805 ;
        RECT 162.355 11.395 162.685 11.725 ;
        RECT 162.355 10.035 162.685 10.365 ;
        RECT 162.355 8.675 162.685 9.005 ;
        RECT 162.355 7.315 162.685 7.645 ;
        RECT 162.355 5.955 162.685 6.285 ;
        RECT 162.355 4.595 162.685 4.925 ;
        RECT 162.355 3.235 162.685 3.565 ;
        RECT 162.355 1.875 162.685 2.205 ;
        RECT 162.355 0.515 162.685 0.845 ;
        RECT 162.36 -8.32 162.68 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.715 15.475 164.045 15.805 ;
        RECT 163.715 10.035 164.045 10.365 ;
        RECT 163.715 8.675 164.045 9.005 ;
        RECT 163.715 7.315 164.045 7.645 ;
        RECT 163.715 5.955 164.045 6.285 ;
        RECT 163.715 4.595 164.045 4.925 ;
        RECT 163.715 3.235 164.045 3.565 ;
        RECT 163.715 1.875 164.045 2.205 ;
        RECT 163.715 0.515 164.045 0.845 ;
        RECT 163.72 -8.32 164.04 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.075 15.475 165.405 15.805 ;
        RECT 165.075 10.035 165.405 10.365 ;
        RECT 165.075 8.675 165.405 9.005 ;
        RECT 165.075 7.315 165.405 7.645 ;
        RECT 165.075 5.955 165.405 6.285 ;
        RECT 165.075 4.595 165.405 4.925 ;
        RECT 165.075 3.235 165.405 3.565 ;
        RECT 165.075 1.875 165.405 2.205 ;
        RECT 165.075 0.515 165.405 0.845 ;
        RECT 165.08 -8.32 165.4 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.435 15.475 166.765 15.805 ;
        RECT 166.435 10.035 166.765 10.365 ;
        RECT 166.435 8.675 166.765 9.005 ;
        RECT 166.435 7.315 166.765 7.645 ;
        RECT 166.435 5.955 166.765 6.285 ;
        RECT 166.435 4.595 166.765 4.925 ;
        RECT 166.435 3.235 166.765 3.565 ;
        RECT 166.435 1.875 166.765 2.205 ;
        RECT 166.435 0.515 166.765 0.845 ;
        RECT 166.44 -8.32 166.76 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.795 15.475 168.125 15.805 ;
        RECT 167.795 10.035 168.125 10.365 ;
        RECT 167.795 8.675 168.125 9.005 ;
        RECT 167.795 7.315 168.125 7.645 ;
        RECT 167.795 5.955 168.125 6.285 ;
        RECT 167.795 4.595 168.125 4.925 ;
        RECT 167.795 3.235 168.125 3.565 ;
        RECT 167.795 1.875 168.125 2.205 ;
        RECT 167.795 0.515 168.125 0.845 ;
        RECT 167.8 -8.32 168.12 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.155 15.475 169.485 15.805 ;
        RECT 169.155 10.035 169.485 10.365 ;
        RECT 169.155 8.675 169.485 9.005 ;
        RECT 169.155 7.315 169.485 7.645 ;
        RECT 169.155 5.955 169.485 6.285 ;
        RECT 169.155 4.595 169.485 4.925 ;
        RECT 169.155 3.235 169.485 3.565 ;
        RECT 169.155 1.875 169.485 2.205 ;
        RECT 169.155 0.515 169.485 0.845 ;
        RECT 169.16 -8.32 169.48 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.515 15.475 170.845 15.805 ;
        RECT 170.515 10.035 170.845 10.365 ;
        RECT 170.515 8.675 170.845 9.005 ;
        RECT 170.515 7.315 170.845 7.645 ;
        RECT 170.515 5.955 170.845 6.285 ;
        RECT 170.515 4.595 170.845 4.925 ;
        RECT 170.515 3.235 170.845 3.565 ;
        RECT 170.515 1.875 170.845 2.205 ;
        RECT 170.515 0.515 170.845 0.845 ;
        RECT 170.52 -8.32 170.84 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.875 15.475 172.205 15.805 ;
        RECT 171.875 11.395 172.205 11.725 ;
        RECT 171.875 10.035 172.205 10.365 ;
        RECT 171.875 8.675 172.205 9.005 ;
        RECT 171.875 7.315 172.205 7.645 ;
        RECT 171.875 5.955 172.205 6.285 ;
        RECT 171.875 4.595 172.205 4.925 ;
        RECT 171.875 3.235 172.205 3.565 ;
        RECT 171.875 1.875 172.205 2.205 ;
        RECT 171.875 0.515 172.205 0.845 ;
        RECT 171.88 -8.32 172.2 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.235 15.475 173.565 15.805 ;
        RECT 173.235 11.395 173.565 11.725 ;
        RECT 173.235 10.035 173.565 10.365 ;
        RECT 173.235 8.675 173.565 9.005 ;
        RECT 173.235 7.315 173.565 7.645 ;
        RECT 173.235 5.955 173.565 6.285 ;
        RECT 173.235 4.595 173.565 4.925 ;
        RECT 173.235 3.235 173.565 3.565 ;
        RECT 173.235 1.875 173.565 2.205 ;
        RECT 173.235 0.515 173.565 0.845 ;
        RECT 173.24 -8.32 173.56 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 174.595 15.475 174.925 15.805 ;
        RECT 174.595 11.395 174.925 11.725 ;
        RECT 174.595 10.035 174.925 10.365 ;
        RECT 174.595 8.675 174.925 9.005 ;
        RECT 174.595 7.315 174.925 7.645 ;
        RECT 174.595 5.955 174.925 6.285 ;
        RECT 174.595 4.595 174.925 4.925 ;
        RECT 174.595 3.235 174.925 3.565 ;
        RECT 174.595 1.875 174.925 2.205 ;
        RECT 174.595 0.515 174.925 0.845 ;
        RECT 174.6 -8.32 174.92 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.955 15.475 176.285 15.805 ;
        RECT 175.955 10.035 176.285 10.365 ;
        RECT 175.955 8.675 176.285 9.005 ;
        RECT 175.955 7.315 176.285 7.645 ;
        RECT 175.955 5.955 176.285 6.285 ;
        RECT 175.955 4.595 176.285 4.925 ;
        RECT 175.955 3.235 176.285 3.565 ;
        RECT 175.955 1.875 176.285 2.205 ;
        RECT 175.955 0.515 176.285 0.845 ;
        RECT 175.96 -8.32 176.28 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.315 15.475 177.645 15.805 ;
        RECT 177.315 10.035 177.645 10.365 ;
        RECT 177.315 8.675 177.645 9.005 ;
        RECT 177.315 7.315 177.645 7.645 ;
        RECT 177.315 5.955 177.645 6.285 ;
        RECT 177.315 4.595 177.645 4.925 ;
        RECT 177.315 3.235 177.645 3.565 ;
        RECT 177.315 1.875 177.645 2.205 ;
        RECT 177.315 0.515 177.645 0.845 ;
        RECT 177.32 -8.32 177.64 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 178.675 15.475 179.005 15.805 ;
        RECT 178.675 10.035 179.005 10.365 ;
        RECT 178.675 8.675 179.005 9.005 ;
        RECT 178.675 7.315 179.005 7.645 ;
        RECT 178.675 5.955 179.005 6.285 ;
        RECT 178.675 4.595 179.005 4.925 ;
        RECT 178.675 3.235 179.005 3.565 ;
        RECT 178.675 1.875 179.005 2.205 ;
        RECT 178.675 0.515 179.005 0.845 ;
        RECT 178.68 -8.32 179 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.035 15.475 180.365 15.805 ;
        RECT 180.035 10.035 180.365 10.365 ;
        RECT 180.035 8.675 180.365 9.005 ;
        RECT 180.035 7.315 180.365 7.645 ;
        RECT 180.035 5.955 180.365 6.285 ;
        RECT 180.035 4.595 180.365 4.925 ;
        RECT 180.035 3.235 180.365 3.565 ;
        RECT 180.035 1.875 180.365 2.205 ;
        RECT 180.035 0.515 180.365 0.845 ;
        RECT 180.04 -8.32 180.36 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 181.395 15.475 181.725 15.805 ;
        RECT 181.395 10.035 181.725 10.365 ;
        RECT 181.395 8.675 181.725 9.005 ;
        RECT 181.395 7.315 181.725 7.645 ;
        RECT 181.395 5.955 181.725 6.285 ;
        RECT 181.395 4.595 181.725 4.925 ;
        RECT 181.395 3.235 181.725 3.565 ;
        RECT 181.395 1.875 181.725 2.205 ;
        RECT 181.395 0.515 181.725 0.845 ;
        RECT 181.4 -8.32 181.72 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.755 15.475 183.085 15.805 ;
        RECT 182.755 10.035 183.085 10.365 ;
        RECT 182.755 8.675 183.085 9.005 ;
        RECT 182.755 7.315 183.085 7.645 ;
        RECT 182.755 5.955 183.085 6.285 ;
        RECT 182.755 4.595 183.085 4.925 ;
        RECT 182.755 3.235 183.085 3.565 ;
        RECT 182.755 1.875 183.085 2.205 ;
        RECT 182.755 0.515 183.085 0.845 ;
        RECT 182.76 -8.32 183.08 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.115 15.475 184.445 15.805 ;
        RECT 184.115 11.395 184.445 11.725 ;
        RECT 184.115 10.035 184.445 10.365 ;
        RECT 184.115 8.675 184.445 9.005 ;
        RECT 184.115 7.315 184.445 7.645 ;
        RECT 184.115 5.955 184.445 6.285 ;
        RECT 184.115 4.595 184.445 4.925 ;
        RECT 184.115 3.235 184.445 3.565 ;
        RECT 184.115 1.875 184.445 2.205 ;
        RECT 184.115 0.515 184.445 0.845 ;
        RECT 184.12 -8.32 184.44 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 185.475 15.475 185.805 15.805 ;
        RECT 185.475 11.395 185.805 11.725 ;
        RECT 185.475 10.035 185.805 10.365 ;
        RECT 185.475 8.675 185.805 9.005 ;
        RECT 185.475 7.315 185.805 7.645 ;
        RECT 185.475 5.955 185.805 6.285 ;
        RECT 185.475 4.595 185.805 4.925 ;
        RECT 185.475 3.235 185.805 3.565 ;
        RECT 185.475 1.875 185.805 2.205 ;
        RECT 185.475 0.515 185.805 0.845 ;
        RECT 185.48 -8.32 185.8 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.835 15.475 187.165 15.805 ;
        RECT 186.835 11.395 187.165 11.725 ;
        RECT 186.835 10.035 187.165 10.365 ;
        RECT 186.835 8.675 187.165 9.005 ;
        RECT 186.835 7.315 187.165 7.645 ;
        RECT 186.835 5.955 187.165 6.285 ;
        RECT 186.835 4.595 187.165 4.925 ;
        RECT 186.835 3.235 187.165 3.565 ;
        RECT 186.835 1.875 187.165 2.205 ;
        RECT 186.835 0.515 187.165 0.845 ;
        RECT 186.84 -8.32 187.16 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.195 15.475 188.525 15.805 ;
        RECT 188.195 10.035 188.525 10.365 ;
        RECT 188.195 8.675 188.525 9.005 ;
        RECT 188.195 7.315 188.525 7.645 ;
        RECT 188.195 5.955 188.525 6.285 ;
        RECT 188.195 4.595 188.525 4.925 ;
        RECT 188.195 3.235 188.525 3.565 ;
        RECT 188.195 1.875 188.525 2.205 ;
        RECT 188.195 0.515 188.525 0.845 ;
        RECT 188.2 -8.32 188.52 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.555 15.475 189.885 15.805 ;
        RECT 189.555 10.035 189.885 10.365 ;
        RECT 189.555 8.675 189.885 9.005 ;
        RECT 189.555 7.315 189.885 7.645 ;
        RECT 189.555 5.955 189.885 6.285 ;
        RECT 189.555 4.595 189.885 4.925 ;
        RECT 189.555 3.235 189.885 3.565 ;
        RECT 189.555 1.875 189.885 2.205 ;
        RECT 189.555 0.515 189.885 0.845 ;
        RECT 189.56 -8.32 189.88 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.915 15.475 191.245 15.805 ;
        RECT 190.915 10.035 191.245 10.365 ;
        RECT 190.915 8.675 191.245 9.005 ;
        RECT 190.915 7.315 191.245 7.645 ;
        RECT 190.915 5.955 191.245 6.285 ;
        RECT 190.915 4.595 191.245 4.925 ;
        RECT 190.915 3.235 191.245 3.565 ;
        RECT 190.915 1.875 191.245 2.205 ;
        RECT 190.915 0.515 191.245 0.845 ;
        RECT 190.92 -8.32 191.24 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.275 15.475 192.605 15.805 ;
        RECT 192.275 10.035 192.605 10.365 ;
        RECT 192.275 8.675 192.605 9.005 ;
        RECT 192.275 7.315 192.605 7.645 ;
        RECT 192.275 5.955 192.605 6.285 ;
        RECT 192.275 4.595 192.605 4.925 ;
        RECT 192.275 3.235 192.605 3.565 ;
        RECT 192.275 1.875 192.605 2.205 ;
        RECT 192.275 0.515 192.605 0.845 ;
        RECT 192.28 -8.32 192.6 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 193.635 15.475 193.965 15.805 ;
        RECT 193.635 10.035 193.965 10.365 ;
        RECT 193.635 8.675 193.965 9.005 ;
        RECT 193.635 7.315 193.965 7.645 ;
        RECT 193.635 5.955 193.965 6.285 ;
        RECT 193.635 4.595 193.965 4.925 ;
        RECT 193.635 3.235 193.965 3.565 ;
        RECT 193.635 1.875 193.965 2.205 ;
        RECT 193.635 0.515 193.965 0.845 ;
        RECT 193.64 -8.32 193.96 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.995 15.475 195.325 15.805 ;
        RECT 194.995 11.395 195.325 11.725 ;
        RECT 194.995 10.035 195.325 10.365 ;
        RECT 194.995 8.675 195.325 9.005 ;
        RECT 194.995 7.315 195.325 7.645 ;
        RECT 194.995 5.955 195.325 6.285 ;
        RECT 194.995 4.595 195.325 4.925 ;
        RECT 194.995 3.235 195.325 3.565 ;
        RECT 194.995 1.875 195.325 2.205 ;
        RECT 194.995 0.515 195.325 0.845 ;
        RECT 195 -8.32 195.32 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 196.355 15.475 196.685 15.805 ;
        RECT 196.355 11.395 196.685 11.725 ;
        RECT 196.355 10.035 196.685 10.365 ;
        RECT 196.355 8.675 196.685 9.005 ;
        RECT 196.355 7.315 196.685 7.645 ;
        RECT 196.355 5.955 196.685 6.285 ;
        RECT 196.355 4.595 196.685 4.925 ;
        RECT 196.355 3.235 196.685 3.565 ;
        RECT 196.355 1.875 196.685 2.205 ;
        RECT 196.355 0.515 196.685 0.845 ;
        RECT 196.36 -8.32 196.68 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.715 15.475 198.045 15.805 ;
        RECT 197.715 11.395 198.045 11.725 ;
        RECT 197.715 10.035 198.045 10.365 ;
        RECT 197.715 8.675 198.045 9.005 ;
        RECT 197.715 7.315 198.045 7.645 ;
        RECT 197.715 5.955 198.045 6.285 ;
        RECT 197.715 4.595 198.045 4.925 ;
        RECT 197.715 3.235 198.045 3.565 ;
        RECT 197.715 1.875 198.045 2.205 ;
        RECT 197.715 0.515 198.045 0.845 ;
        RECT 197.72 -8.32 198.04 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.075 15.475 199.405 15.805 ;
        RECT 199.075 10.035 199.405 10.365 ;
        RECT 199.075 8.675 199.405 9.005 ;
        RECT 199.075 7.315 199.405 7.645 ;
        RECT 199.075 5.955 199.405 6.285 ;
        RECT 199.075 4.595 199.405 4.925 ;
        RECT 199.075 3.235 199.405 3.565 ;
        RECT 199.075 1.875 199.405 2.205 ;
        RECT 199.075 0.515 199.405 0.845 ;
        RECT 199.08 -8.32 199.4 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 200.435 15.475 200.765 15.805 ;
        RECT 200.435 10.035 200.765 10.365 ;
        RECT 200.435 8.675 200.765 9.005 ;
        RECT 200.435 7.315 200.765 7.645 ;
        RECT 200.435 5.955 200.765 6.285 ;
        RECT 200.435 4.595 200.765 4.925 ;
        RECT 200.435 3.235 200.765 3.565 ;
        RECT 200.435 1.875 200.765 2.205 ;
        RECT 200.435 0.515 200.765 0.845 ;
        RECT 200.44 -8.32 200.76 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.795 15.475 202.125 15.805 ;
        RECT 201.795 10.035 202.125 10.365 ;
        RECT 201.795 8.675 202.125 9.005 ;
        RECT 201.795 7.315 202.125 7.645 ;
        RECT 201.795 5.955 202.125 6.285 ;
        RECT 201.795 4.595 202.125 4.925 ;
        RECT 201.795 3.235 202.125 3.565 ;
        RECT 201.795 1.875 202.125 2.205 ;
        RECT 201.795 0.515 202.125 0.845 ;
        RECT 201.8 -8.32 202.12 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.155 15.475 203.485 15.805 ;
        RECT 203.155 10.035 203.485 10.365 ;
        RECT 203.155 8.675 203.485 9.005 ;
        RECT 203.155 7.315 203.485 7.645 ;
        RECT 203.155 5.955 203.485 6.285 ;
        RECT 203.155 4.595 203.485 4.925 ;
        RECT 203.155 3.235 203.485 3.565 ;
        RECT 203.155 1.875 203.485 2.205 ;
        RECT 203.155 0.515 203.485 0.845 ;
        RECT 203.16 -8.32 203.48 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 204.515 15.475 204.845 15.805 ;
        RECT 204.515 10.035 204.845 10.365 ;
        RECT 204.515 8.675 204.845 9.005 ;
        RECT 204.515 7.315 204.845 7.645 ;
        RECT 204.515 5.955 204.845 6.285 ;
        RECT 204.515 4.595 204.845 4.925 ;
        RECT 204.515 3.235 204.845 3.565 ;
        RECT 204.515 1.875 204.845 2.205 ;
        RECT 204.515 0.515 204.845 0.845 ;
        RECT 204.52 -8.32 204.84 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.875 15.475 206.205 15.805 ;
        RECT 205.875 10.035 206.205 10.365 ;
        RECT 205.875 8.675 206.205 9.005 ;
        RECT 205.875 7.315 206.205 7.645 ;
        RECT 205.875 5.955 206.205 6.285 ;
        RECT 205.875 4.595 206.205 4.925 ;
        RECT 205.875 3.235 206.205 3.565 ;
        RECT 205.875 1.875 206.205 2.205 ;
        RECT 205.875 0.515 206.205 0.845 ;
        RECT 205.88 -8.32 206.2 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.235 15.475 207.565 15.805 ;
        RECT 207.235 11.395 207.565 11.725 ;
        RECT 207.235 10.035 207.565 10.365 ;
        RECT 207.235 8.675 207.565 9.005 ;
        RECT 207.235 7.315 207.565 7.645 ;
        RECT 207.235 5.955 207.565 6.285 ;
        RECT 207.235 4.595 207.565 4.925 ;
        RECT 207.235 3.235 207.565 3.565 ;
        RECT 207.235 1.875 207.565 2.205 ;
        RECT 207.235 0.515 207.565 0.845 ;
        RECT 207.24 -8.32 207.56 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 208.595 15.475 208.925 15.805 ;
        RECT 208.595 11.395 208.925 11.725 ;
        RECT 208.595 10.035 208.925 10.365 ;
        RECT 208.595 8.675 208.925 9.005 ;
        RECT 208.595 7.315 208.925 7.645 ;
        RECT 208.595 5.955 208.925 6.285 ;
        RECT 208.595 4.595 208.925 4.925 ;
        RECT 208.595 3.235 208.925 3.565 ;
        RECT 208.595 1.875 208.925 2.205 ;
        RECT 208.595 0.515 208.925 0.845 ;
        RECT 208.6 -8.32 208.92 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.955 15.475 210.285 15.805 ;
        RECT 209.955 11.395 210.285 11.725 ;
        RECT 209.955 10.035 210.285 10.365 ;
        RECT 209.955 8.675 210.285 9.005 ;
        RECT 209.955 7.315 210.285 7.645 ;
        RECT 209.955 5.955 210.285 6.285 ;
        RECT 209.955 4.595 210.285 4.925 ;
        RECT 209.955 3.235 210.285 3.565 ;
        RECT 209.955 1.875 210.285 2.205 ;
        RECT 209.955 0.515 210.285 0.845 ;
        RECT 209.96 -8.32 210.28 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 211.315 15.475 211.645 15.805 ;
        RECT 211.315 10.035 211.645 10.365 ;
        RECT 211.315 8.675 211.645 9.005 ;
        RECT 211.315 7.315 211.645 7.645 ;
        RECT 211.315 5.955 211.645 6.285 ;
        RECT 211.315 4.595 211.645 4.925 ;
        RECT 211.315 3.235 211.645 3.565 ;
        RECT 211.315 1.875 211.645 2.205 ;
        RECT 211.315 0.515 211.645 0.845 ;
        RECT 211.32 -8.32 211.64 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 212.675 15.475 213.005 15.805 ;
        RECT 212.675 10.035 213.005 10.365 ;
        RECT 212.675 8.675 213.005 9.005 ;
        RECT 212.675 7.315 213.005 7.645 ;
        RECT 212.675 5.955 213.005 6.285 ;
        RECT 212.675 4.595 213.005 4.925 ;
        RECT 212.675 3.235 213.005 3.565 ;
        RECT 212.675 1.875 213.005 2.205 ;
        RECT 212.675 0.515 213.005 0.845 ;
        RECT 212.68 -8.32 213 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.035 15.475 214.365 15.805 ;
        RECT 214.035 10.035 214.365 10.365 ;
        RECT 214.035 8.675 214.365 9.005 ;
        RECT 214.035 7.315 214.365 7.645 ;
        RECT 214.035 5.955 214.365 6.285 ;
        RECT 214.035 4.595 214.365 4.925 ;
        RECT 214.035 3.235 214.365 3.565 ;
        RECT 214.035 1.875 214.365 2.205 ;
        RECT 214.035 0.515 214.365 0.845 ;
        RECT 214.04 -8.32 214.36 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 215.395 15.475 215.725 15.805 ;
        RECT 215.395 10.035 215.725 10.365 ;
        RECT 215.395 8.675 215.725 9.005 ;
        RECT 215.395 7.315 215.725 7.645 ;
        RECT 215.395 5.955 215.725 6.285 ;
        RECT 215.395 4.595 215.725 4.925 ;
        RECT 215.395 3.235 215.725 3.565 ;
        RECT 215.395 1.875 215.725 2.205 ;
        RECT 215.395 0.515 215.725 0.845 ;
        RECT 215.4 -8.32 215.72 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.755 15.475 217.085 15.805 ;
        RECT 216.755 10.035 217.085 10.365 ;
        RECT 216.755 8.675 217.085 9.005 ;
        RECT 216.755 7.315 217.085 7.645 ;
        RECT 216.755 5.955 217.085 6.285 ;
        RECT 216.755 4.595 217.085 4.925 ;
        RECT 216.755 3.235 217.085 3.565 ;
        RECT 216.755 1.875 217.085 2.205 ;
        RECT 216.755 0.515 217.085 0.845 ;
        RECT 216.76 -8.32 217.08 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.115 15.475 218.445 15.805 ;
        RECT 218.115 10.035 218.445 10.365 ;
        RECT 218.115 8.675 218.445 9.005 ;
        RECT 218.115 7.315 218.445 7.645 ;
        RECT 218.115 5.955 218.445 6.285 ;
        RECT 218.115 4.595 218.445 4.925 ;
        RECT 218.115 3.235 218.445 3.565 ;
        RECT 218.115 1.875 218.445 2.205 ;
        RECT 218.115 0.515 218.445 0.845 ;
        RECT 218.12 -8.32 218.44 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 219.475 15.475 219.805 15.805 ;
        RECT 219.475 11.395 219.805 11.725 ;
        RECT 219.475 10.035 219.805 10.365 ;
        RECT 219.475 8.675 219.805 9.005 ;
        RECT 219.475 7.315 219.805 7.645 ;
        RECT 219.475 5.955 219.805 6.285 ;
        RECT 219.475 4.595 219.805 4.925 ;
        RECT 219.475 3.235 219.805 3.565 ;
        RECT 219.475 1.875 219.805 2.205 ;
        RECT 219.475 0.515 219.805 0.845 ;
        RECT 219.48 -8.32 219.8 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.835 15.475 221.165 15.805 ;
        RECT 220.835 11.395 221.165 11.725 ;
        RECT 220.835 10.035 221.165 10.365 ;
        RECT 220.835 8.675 221.165 9.005 ;
        RECT 220.835 7.315 221.165 7.645 ;
        RECT 220.835 5.955 221.165 6.285 ;
        RECT 220.835 4.595 221.165 4.925 ;
        RECT 220.835 3.235 221.165 3.565 ;
        RECT 220.835 1.875 221.165 2.205 ;
        RECT 220.835 0.515 221.165 0.845 ;
        RECT 220.84 -8.32 221.16 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.195 15.475 222.525 15.805 ;
        RECT 222.195 11.395 222.525 11.725 ;
        RECT 222.195 10.035 222.525 10.365 ;
        RECT 222.195 8.675 222.525 9.005 ;
        RECT 222.195 7.315 222.525 7.645 ;
        RECT 222.195 5.955 222.525 6.285 ;
        RECT 222.195 4.595 222.525 4.925 ;
        RECT 222.195 3.235 222.525 3.565 ;
        RECT 222.195 1.875 222.525 2.205 ;
        RECT 222.195 0.515 222.525 0.845 ;
        RECT 222.2 -8.32 222.52 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 223.555 15.475 223.885 15.805 ;
        RECT 223.555 10.035 223.885 10.365 ;
        RECT 223.555 8.675 223.885 9.005 ;
        RECT 223.555 7.315 223.885 7.645 ;
        RECT 223.555 5.955 223.885 6.285 ;
        RECT 223.555 4.595 223.885 4.925 ;
        RECT 223.555 3.235 223.885 3.565 ;
        RECT 223.555 1.875 223.885 2.205 ;
        RECT 223.555 0.515 223.885 0.845 ;
        RECT 223.56 -8.32 223.88 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 224.915 15.475 225.245 15.805 ;
        RECT 224.915 10.035 225.245 10.365 ;
        RECT 224.915 8.675 225.245 9.005 ;
        RECT 224.915 7.315 225.245 7.645 ;
        RECT 224.915 5.955 225.245 6.285 ;
        RECT 224.915 4.595 225.245 4.925 ;
        RECT 224.915 3.235 225.245 3.565 ;
        RECT 224.915 1.875 225.245 2.205 ;
        RECT 224.915 0.515 225.245 0.845 ;
        RECT 224.92 -8.32 225.24 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.275 15.475 226.605 15.805 ;
        RECT 226.275 10.035 226.605 10.365 ;
        RECT 226.275 8.675 226.605 9.005 ;
        RECT 226.275 7.315 226.605 7.645 ;
        RECT 226.275 5.955 226.605 6.285 ;
        RECT 226.275 4.595 226.605 4.925 ;
        RECT 226.275 3.235 226.605 3.565 ;
        RECT 226.275 1.875 226.605 2.205 ;
        RECT 226.275 0.515 226.605 0.845 ;
        RECT 226.28 -8.32 226.6 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 227.635 15.475 227.965 15.805 ;
        RECT 227.635 10.035 227.965 10.365 ;
        RECT 227.635 8.675 227.965 9.005 ;
        RECT 227.635 7.315 227.965 7.645 ;
        RECT 227.635 5.955 227.965 6.285 ;
        RECT 227.635 4.595 227.965 4.925 ;
        RECT 227.635 3.235 227.965 3.565 ;
        RECT 227.635 1.875 227.965 2.205 ;
        RECT 227.635 0.515 227.965 0.845 ;
        RECT 227.64 -8.32 227.96 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.995 15.475 229.325 15.805 ;
        RECT 228.995 10.035 229.325 10.365 ;
        RECT 228.995 8.675 229.325 9.005 ;
        RECT 228.995 7.315 229.325 7.645 ;
        RECT 228.995 5.955 229.325 6.285 ;
        RECT 228.995 4.595 229.325 4.925 ;
        RECT 228.995 3.235 229.325 3.565 ;
        RECT 228.995 1.875 229.325 2.205 ;
        RECT 228.995 0.515 229.325 0.845 ;
        RECT 229 -8.32 229.32 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 230.355 15.475 230.685 15.805 ;
        RECT 230.355 10.035 230.685 10.365 ;
        RECT 230.355 8.675 230.685 9.005 ;
        RECT 230.355 7.315 230.685 7.645 ;
        RECT 230.355 5.955 230.685 6.285 ;
        RECT 230.355 4.595 230.685 4.925 ;
        RECT 230.355 3.235 230.685 3.565 ;
        RECT 230.355 1.875 230.685 2.205 ;
        RECT 230.355 0.515 230.685 0.845 ;
        RECT 230.36 -8.32 230.68 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 231.715 15.475 232.045 15.805 ;
        RECT 231.715 11.395 232.045 11.725 ;
        RECT 231.715 10.035 232.045 10.365 ;
        RECT 231.715 8.675 232.045 9.005 ;
        RECT 231.715 7.315 232.045 7.645 ;
        RECT 231.715 5.955 232.045 6.285 ;
        RECT 231.715 4.595 232.045 4.925 ;
        RECT 231.715 3.235 232.045 3.565 ;
        RECT 231.715 1.875 232.045 2.205 ;
        RECT 231.715 0.515 232.045 0.845 ;
        RECT 231.72 -8.32 232.04 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.075 15.475 233.405 15.805 ;
        RECT 233.075 11.395 233.405 11.725 ;
        RECT 233.075 10.035 233.405 10.365 ;
        RECT 233.075 8.675 233.405 9.005 ;
        RECT 233.075 7.315 233.405 7.645 ;
        RECT 233.075 5.955 233.405 6.285 ;
        RECT 233.075 4.595 233.405 4.925 ;
        RECT 233.075 3.235 233.405 3.565 ;
        RECT 233.075 1.875 233.405 2.205 ;
        RECT 233.075 0.515 233.405 0.845 ;
        RECT 233.08 -8.32 233.4 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 234.435 15.475 234.765 15.805 ;
        RECT 234.435 11.395 234.765 11.725 ;
        RECT 234.435 10.035 234.765 10.365 ;
        RECT 234.435 8.675 234.765 9.005 ;
        RECT 234.435 7.315 234.765 7.645 ;
        RECT 234.435 5.955 234.765 6.285 ;
        RECT 234.435 4.595 234.765 4.925 ;
        RECT 234.435 3.235 234.765 3.565 ;
        RECT 234.435 1.875 234.765 2.205 ;
        RECT 234.435 0.515 234.765 0.845 ;
        RECT 234.44 -8.32 234.76 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 235.795 15.475 236.125 15.805 ;
        RECT 235.795 10.035 236.125 10.365 ;
        RECT 235.795 8.675 236.125 9.005 ;
        RECT 235.795 7.315 236.125 7.645 ;
        RECT 235.795 5.955 236.125 6.285 ;
        RECT 235.795 4.595 236.125 4.925 ;
        RECT 235.795 3.235 236.125 3.565 ;
        RECT 235.795 1.875 236.125 2.205 ;
        RECT 235.795 0.515 236.125 0.845 ;
        RECT 235.8 -8.32 236.12 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 237.155 15.475 237.485 15.805 ;
        RECT 237.155 10.035 237.485 10.365 ;
        RECT 237.155 8.675 237.485 9.005 ;
        RECT 237.155 7.315 237.485 7.645 ;
        RECT 237.155 5.955 237.485 6.285 ;
        RECT 237.155 4.595 237.485 4.925 ;
        RECT 237.155 3.235 237.485 3.565 ;
        RECT 237.155 1.875 237.485 2.205 ;
        RECT 237.155 0.515 237.485 0.845 ;
        RECT 237.16 -8.32 237.48 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 238.515 15.475 238.845 15.805 ;
        RECT 238.515 10.035 238.845 10.365 ;
        RECT 238.515 8.675 238.845 9.005 ;
        RECT 238.515 7.315 238.845 7.645 ;
        RECT 238.515 5.955 238.845 6.285 ;
        RECT 238.515 4.595 238.845 4.925 ;
        RECT 238.515 3.235 238.845 3.565 ;
        RECT 238.515 1.875 238.845 2.205 ;
        RECT 238.515 0.515 238.845 0.845 ;
        RECT 238.52 -8.32 238.84 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.875 15.475 240.205 15.805 ;
        RECT 239.875 10.035 240.205 10.365 ;
        RECT 239.875 8.675 240.205 9.005 ;
        RECT 239.875 7.315 240.205 7.645 ;
        RECT 239.875 5.955 240.205 6.285 ;
        RECT 239.875 4.595 240.205 4.925 ;
        RECT 239.875 3.235 240.205 3.565 ;
        RECT 239.875 1.875 240.205 2.205 ;
        RECT 239.875 0.515 240.205 0.845 ;
        RECT 239.88 -8.32 240.2 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 241.235 15.475 241.565 15.805 ;
        RECT 241.235 10.035 241.565 10.365 ;
        RECT 241.235 8.675 241.565 9.005 ;
        RECT 241.235 7.315 241.565 7.645 ;
        RECT 241.235 5.955 241.565 6.285 ;
        RECT 241.235 4.595 241.565 4.925 ;
        RECT 241.235 3.235 241.565 3.565 ;
        RECT 241.235 1.875 241.565 2.205 ;
        RECT 241.235 0.515 241.565 0.845 ;
        RECT 241.24 -8.32 241.56 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 242.595 15.475 242.925 15.805 ;
        RECT 242.595 10.035 242.925 10.365 ;
        RECT 242.595 8.675 242.925 9.005 ;
        RECT 242.595 7.315 242.925 7.645 ;
        RECT 242.595 5.955 242.925 6.285 ;
        RECT 242.595 4.595 242.925 4.925 ;
        RECT 242.595 3.235 242.925 3.565 ;
        RECT 242.595 1.875 242.925 2.205 ;
        RECT 242.595 0.515 242.925 0.845 ;
        RECT 242.6 -8.32 242.92 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 243.955 15.475 244.285 15.805 ;
        RECT 243.955 11.395 244.285 11.725 ;
        RECT 243.955 10.035 244.285 10.365 ;
        RECT 243.955 8.675 244.285 9.005 ;
        RECT 243.955 7.315 244.285 7.645 ;
        RECT 243.955 5.955 244.285 6.285 ;
        RECT 243.955 4.595 244.285 4.925 ;
        RECT 243.955 3.235 244.285 3.565 ;
        RECT 243.955 1.875 244.285 2.205 ;
        RECT 243.955 0.515 244.285 0.845 ;
        RECT 243.96 -8.32 244.28 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 245.315 0.515 245.645 0.845 ;
        RECT 245.32 -8.32 245.64 15.805 ;
        RECT 245.315 15.475 245.645 15.805 ;
        RECT 245.315 11.395 245.645 11.725 ;
        RECT 245.315 10.035 245.645 10.365 ;
        RECT 245.315 8.675 245.645 9.005 ;
        RECT 245.315 7.315 245.645 7.645 ;
        RECT 245.315 5.955 245.645 6.285 ;
        RECT 245.315 4.595 245.645 4.925 ;
        RECT 245.315 3.235 245.645 3.565 ;
        RECT 245.315 1.875 245.645 2.205 ;
    END
    PORT
      LAYER met3 ;
        RECT -2.205 15.475 -1.875 15.805 ;
        RECT -2.205 14.115 -1.875 14.445 ;
        RECT -2.205 12.755 -1.875 13.085 ;
        RECT -2.205 11.395 -1.875 11.725 ;
        RECT -2.205 10.035 -1.875 10.365 ;
        RECT -2.205 8.675 -1.875 9.005 ;
        RECT -2.205 7.315 -1.875 7.645 ;
        RECT -2.205 5.955 -1.875 6.285 ;
        RECT -2.205 4.595 -1.875 4.925 ;
        RECT -2.205 3.235 -1.875 3.565 ;
        RECT -2.205 1.875 -1.875 2.205 ;
        RECT -2.205 0.515 -1.875 0.845 ;
        RECT -2.2 -8.32 -1.88 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.845 15.475 -0.515 15.805 ;
        RECT -0.845 14.115 -0.515 14.445 ;
        RECT -0.845 12.755 -0.515 13.085 ;
        RECT -0.845 11.395 -0.515 11.725 ;
        RECT -0.845 10.035 -0.515 10.365 ;
        RECT -0.845 8.675 -0.515 9.005 ;
        RECT -0.845 7.315 -0.515 7.645 ;
        RECT -0.845 5.955 -0.515 6.285 ;
        RECT -0.845 4.595 -0.515 4.925 ;
        RECT -0.845 3.235 -0.515 3.565 ;
        RECT -0.845 1.875 -0.515 2.205 ;
        RECT -0.845 0.515 -0.515 0.845 ;
        RECT -0.84 -8.32 -0.52 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.515 15.475 0.845 15.805 ;
        RECT 0.515 12.755 0.845 13.085 ;
        RECT 0.515 11.395 0.845 11.725 ;
        RECT 0.515 10.035 0.845 10.365 ;
        RECT 0.515 8.675 0.845 9.005 ;
        RECT 0.515 7.315 0.845 7.645 ;
        RECT 0.515 5.955 0.845 6.285 ;
        RECT 0.515 4.595 0.845 4.925 ;
        RECT 0.515 3.235 0.845 3.565 ;
        RECT 0.515 1.875 0.845 2.205 ;
        RECT 0.515 0.515 0.845 0.845 ;
        RECT 0.52 -8.32 0.84 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.875 15.475 2.205 15.805 ;
        RECT 1.875 11.395 2.205 11.725 ;
        RECT 1.875 10.035 2.205 10.365 ;
        RECT 1.875 8.675 2.205 9.005 ;
        RECT 1.875 7.315 2.205 7.645 ;
        RECT 1.875 5.955 2.205 6.285 ;
        RECT 1.875 4.595 2.205 4.925 ;
        RECT 1.875 3.235 2.205 3.565 ;
        RECT 1.875 1.875 2.205 2.205 ;
        RECT 1.875 0.515 2.205 0.845 ;
        RECT 1.88 -8.32 2.2 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.235 15.475 3.565 15.805 ;
        RECT 3.235 11.395 3.565 11.725 ;
        RECT 3.235 10.035 3.565 10.365 ;
        RECT 3.235 8.675 3.565 9.005 ;
        RECT 3.235 7.315 3.565 7.645 ;
        RECT 3.235 5.955 3.565 6.285 ;
        RECT 3.235 4.595 3.565 4.925 ;
        RECT 3.235 3.235 3.565 3.565 ;
        RECT 3.235 1.875 3.565 2.205 ;
        RECT 3.235 0.515 3.565 0.845 ;
        RECT 3.24 -8.32 3.56 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.595 15.475 4.925 15.805 ;
        RECT 4.595 11.395 4.925 11.725 ;
        RECT 4.595 10.035 4.925 10.365 ;
        RECT 4.595 8.675 4.925 9.005 ;
        RECT 4.595 7.315 4.925 7.645 ;
        RECT 4.595 5.955 4.925 6.285 ;
        RECT 4.595 4.595 4.925 4.925 ;
        RECT 4.595 3.235 4.925 3.565 ;
        RECT 4.595 1.875 4.925 2.205 ;
        RECT 4.595 0.515 4.925 0.845 ;
        RECT 4.6 -8.32 4.92 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.955 15.475 6.285 15.805 ;
        RECT 5.955 11.395 6.285 11.725 ;
        RECT 5.955 10.035 6.285 10.365 ;
        RECT 5.955 8.675 6.285 9.005 ;
        RECT 5.955 7.315 6.285 7.645 ;
        RECT 5.955 5.955 6.285 6.285 ;
        RECT 5.955 4.595 6.285 4.925 ;
        RECT 5.955 3.235 6.285 3.565 ;
        RECT 5.955 1.875 6.285 2.205 ;
        RECT 5.955 0.515 6.285 0.845 ;
        RECT 5.96 -8.32 6.28 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.315 15.475 7.645 15.805 ;
        RECT 7.315 10.035 7.645 10.365 ;
        RECT 7.315 8.675 7.645 9.005 ;
        RECT 7.315 7.315 7.645 7.645 ;
        RECT 7.315 5.955 7.645 6.285 ;
        RECT 7.315 4.595 7.645 4.925 ;
        RECT 7.315 3.235 7.645 3.565 ;
        RECT 7.315 1.875 7.645 2.205 ;
        RECT 7.315 0.515 7.645 0.845 ;
        RECT 7.32 -8.32 7.64 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.675 15.475 9.005 15.805 ;
        RECT 8.675 10.035 9.005 10.365 ;
        RECT 8.675 8.675 9.005 9.005 ;
        RECT 8.675 7.315 9.005 7.645 ;
        RECT 8.675 5.955 9.005 6.285 ;
        RECT 8.675 4.595 9.005 4.925 ;
        RECT 8.675 3.235 9.005 3.565 ;
        RECT 8.675 1.875 9.005 2.205 ;
        RECT 8.675 0.515 9.005 0.845 ;
        RECT 8.68 -8.32 9 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.035 15.475 10.365 15.805 ;
        RECT 10.035 10.035 10.365 10.365 ;
        RECT 10.035 8.675 10.365 9.005 ;
        RECT 10.035 7.315 10.365 7.645 ;
        RECT 10.035 5.955 10.365 6.285 ;
        RECT 10.035 4.595 10.365 4.925 ;
        RECT 10.035 3.235 10.365 3.565 ;
        RECT 10.035 1.875 10.365 2.205 ;
        RECT 10.035 0.515 10.365 0.845 ;
        RECT 10.04 -8.32 10.36 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.395 15.475 11.725 15.805 ;
        RECT 11.395 10.035 11.725 10.365 ;
        RECT 11.395 8.675 11.725 9.005 ;
        RECT 11.395 7.315 11.725 7.645 ;
        RECT 11.395 5.955 11.725 6.285 ;
        RECT 11.395 4.595 11.725 4.925 ;
        RECT 11.395 3.235 11.725 3.565 ;
        RECT 11.395 1.875 11.725 2.205 ;
        RECT 11.395 0.515 11.725 0.845 ;
        RECT 11.4 -8.32 11.72 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.755 15.475 13.085 15.805 ;
        RECT 12.755 10.035 13.085 10.365 ;
        RECT 12.755 8.675 13.085 9.005 ;
        RECT 12.755 7.315 13.085 7.645 ;
        RECT 12.755 5.955 13.085 6.285 ;
        RECT 12.755 4.595 13.085 4.925 ;
        RECT 12.755 3.235 13.085 3.565 ;
        RECT 12.755 1.875 13.085 2.205 ;
        RECT 12.755 0.515 13.085 0.845 ;
        RECT 12.76 -8.32 13.08 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.115 15.475 14.445 15.805 ;
        RECT 14.115 10.035 14.445 10.365 ;
        RECT 14.115 8.675 14.445 9.005 ;
        RECT 14.115 7.315 14.445 7.645 ;
        RECT 14.115 5.955 14.445 6.285 ;
        RECT 14.115 4.595 14.445 4.925 ;
        RECT 14.115 3.235 14.445 3.565 ;
        RECT 14.115 1.875 14.445 2.205 ;
        RECT 14.115 0.515 14.445 0.845 ;
        RECT 14.12 -8.32 14.44 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.475 15.475 15.805 15.805 ;
        RECT 15.475 11.395 15.805 11.725 ;
        RECT 15.475 10.035 15.805 10.365 ;
        RECT 15.475 8.675 15.805 9.005 ;
        RECT 15.475 7.315 15.805 7.645 ;
        RECT 15.475 5.955 15.805 6.285 ;
        RECT 15.475 4.595 15.805 4.925 ;
        RECT 15.475 3.235 15.805 3.565 ;
        RECT 15.475 1.875 15.805 2.205 ;
        RECT 15.475 0.515 15.805 0.845 ;
        RECT 15.48 -8.32 15.8 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.835 15.475 17.165 15.805 ;
        RECT 16.835 11.395 17.165 11.725 ;
        RECT 16.835 10.035 17.165 10.365 ;
        RECT 16.835 8.675 17.165 9.005 ;
        RECT 16.835 7.315 17.165 7.645 ;
        RECT 16.835 5.955 17.165 6.285 ;
        RECT 16.835 4.595 17.165 4.925 ;
        RECT 16.835 3.235 17.165 3.565 ;
        RECT 16.835 1.875 17.165 2.205 ;
        RECT 16.835 0.515 17.165 0.845 ;
        RECT 16.84 -8.32 17.16 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.195 15.475 18.525 15.805 ;
        RECT 18.195 11.395 18.525 11.725 ;
        RECT 18.195 10.035 18.525 10.365 ;
        RECT 18.195 8.675 18.525 9.005 ;
        RECT 18.195 7.315 18.525 7.645 ;
        RECT 18.195 5.955 18.525 6.285 ;
        RECT 18.195 4.595 18.525 4.925 ;
        RECT 18.195 3.235 18.525 3.565 ;
        RECT 18.195 1.875 18.525 2.205 ;
        RECT 18.195 0.515 18.525 0.845 ;
        RECT 18.2 -8.32 18.52 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.555 15.475 19.885 15.805 ;
        RECT 19.555 10.035 19.885 10.365 ;
        RECT 19.555 8.675 19.885 9.005 ;
        RECT 19.555 7.315 19.885 7.645 ;
        RECT 19.555 5.955 19.885 6.285 ;
        RECT 19.555 4.595 19.885 4.925 ;
        RECT 19.555 3.235 19.885 3.565 ;
        RECT 19.555 1.875 19.885 2.205 ;
        RECT 19.555 0.515 19.885 0.845 ;
        RECT 19.56 -8.32 19.88 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.915 15.475 21.245 15.805 ;
        RECT 20.915 10.035 21.245 10.365 ;
        RECT 20.915 8.675 21.245 9.005 ;
        RECT 20.915 7.315 21.245 7.645 ;
        RECT 20.915 5.955 21.245 6.285 ;
        RECT 20.915 4.595 21.245 4.925 ;
        RECT 20.915 3.235 21.245 3.565 ;
        RECT 20.915 1.875 21.245 2.205 ;
        RECT 20.915 0.515 21.245 0.845 ;
        RECT 20.92 -8.32 21.24 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.275 15.475 22.605 15.805 ;
        RECT 22.275 10.035 22.605 10.365 ;
        RECT 22.275 8.675 22.605 9.005 ;
        RECT 22.275 7.315 22.605 7.645 ;
        RECT 22.275 5.955 22.605 6.285 ;
        RECT 22.275 4.595 22.605 4.925 ;
        RECT 22.275 3.235 22.605 3.565 ;
        RECT 22.275 1.875 22.605 2.205 ;
        RECT 22.275 0.515 22.605 0.845 ;
        RECT 22.28 -8.32 22.6 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.635 15.475 23.965 15.805 ;
        RECT 23.635 10.035 23.965 10.365 ;
        RECT 23.635 8.675 23.965 9.005 ;
        RECT 23.635 7.315 23.965 7.645 ;
        RECT 23.635 5.955 23.965 6.285 ;
        RECT 23.635 4.595 23.965 4.925 ;
        RECT 23.635 3.235 23.965 3.565 ;
        RECT 23.635 1.875 23.965 2.205 ;
        RECT 23.635 0.515 23.965 0.845 ;
        RECT 23.64 -8.32 23.96 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.995 15.475 25.325 15.805 ;
        RECT 24.995 10.035 25.325 10.365 ;
        RECT 24.995 8.675 25.325 9.005 ;
        RECT 24.995 7.315 25.325 7.645 ;
        RECT 24.995 5.955 25.325 6.285 ;
        RECT 24.995 4.595 25.325 4.925 ;
        RECT 24.995 3.235 25.325 3.565 ;
        RECT 24.995 1.875 25.325 2.205 ;
        RECT 24.995 0.515 25.325 0.845 ;
        RECT 25 -8.32 25.32 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.355 15.475 26.685 15.805 ;
        RECT 26.355 10.035 26.685 10.365 ;
        RECT 26.355 8.675 26.685 9.005 ;
        RECT 26.355 7.315 26.685 7.645 ;
        RECT 26.355 5.955 26.685 6.285 ;
        RECT 26.355 4.595 26.685 4.925 ;
        RECT 26.355 3.235 26.685 3.565 ;
        RECT 26.355 1.875 26.685 2.205 ;
        RECT 26.355 0.515 26.685 0.845 ;
        RECT 26.36 -8.32 26.68 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.715 15.475 28.045 15.805 ;
        RECT 27.715 11.395 28.045 11.725 ;
        RECT 27.715 10.035 28.045 10.365 ;
        RECT 27.715 8.675 28.045 9.005 ;
        RECT 27.715 7.315 28.045 7.645 ;
        RECT 27.715 5.955 28.045 6.285 ;
        RECT 27.715 4.595 28.045 4.925 ;
        RECT 27.715 3.235 28.045 3.565 ;
        RECT 27.715 1.875 28.045 2.205 ;
        RECT 27.715 0.515 28.045 0.845 ;
        RECT 27.72 -8.32 28.04 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.075 15.475 29.405 15.805 ;
        RECT 29.075 11.395 29.405 11.725 ;
        RECT 29.075 10.035 29.405 10.365 ;
        RECT 29.075 8.675 29.405 9.005 ;
        RECT 29.075 7.315 29.405 7.645 ;
        RECT 29.075 5.955 29.405 6.285 ;
        RECT 29.075 4.595 29.405 4.925 ;
        RECT 29.075 3.235 29.405 3.565 ;
        RECT 29.075 1.875 29.405 2.205 ;
        RECT 29.075 0.515 29.405 0.845 ;
        RECT 29.08 -8.32 29.4 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.435 15.475 30.765 15.805 ;
        RECT 30.435 11.395 30.765 11.725 ;
        RECT 30.435 10.035 30.765 10.365 ;
        RECT 30.435 8.675 30.765 9.005 ;
        RECT 30.435 7.315 30.765 7.645 ;
        RECT 30.435 5.955 30.765 6.285 ;
        RECT 30.435 4.595 30.765 4.925 ;
        RECT 30.435 3.235 30.765 3.565 ;
        RECT 30.435 1.875 30.765 2.205 ;
        RECT 30.435 0.515 30.765 0.845 ;
        RECT 30.44 -8.32 30.76 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.795 15.475 32.125 15.805 ;
        RECT 31.795 10.035 32.125 10.365 ;
        RECT 31.795 8.675 32.125 9.005 ;
        RECT 31.795 7.315 32.125 7.645 ;
        RECT 31.795 5.955 32.125 6.285 ;
        RECT 31.795 4.595 32.125 4.925 ;
        RECT 31.795 3.235 32.125 3.565 ;
        RECT 31.795 1.875 32.125 2.205 ;
        RECT 31.795 0.515 32.125 0.845 ;
        RECT 31.8 -8.32 32.12 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.155 15.475 33.485 15.805 ;
        RECT 33.155 10.035 33.485 10.365 ;
        RECT 33.155 8.675 33.485 9.005 ;
        RECT 33.155 7.315 33.485 7.645 ;
        RECT 33.155 5.955 33.485 6.285 ;
        RECT 33.155 4.595 33.485 4.925 ;
        RECT 33.155 3.235 33.485 3.565 ;
        RECT 33.155 1.875 33.485 2.205 ;
        RECT 33.155 0.515 33.485 0.845 ;
        RECT 33.16 -8.32 33.48 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.515 15.475 34.845 15.805 ;
        RECT 34.515 10.035 34.845 10.365 ;
        RECT 34.515 8.675 34.845 9.005 ;
        RECT 34.515 7.315 34.845 7.645 ;
        RECT 34.515 5.955 34.845 6.285 ;
        RECT 34.515 4.595 34.845 4.925 ;
        RECT 34.515 3.235 34.845 3.565 ;
        RECT 34.515 1.875 34.845 2.205 ;
        RECT 34.515 0.515 34.845 0.845 ;
        RECT 34.52 -8.32 34.84 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.875 15.475 36.205 15.805 ;
        RECT 35.875 10.035 36.205 10.365 ;
        RECT 35.875 8.675 36.205 9.005 ;
        RECT 35.875 7.315 36.205 7.645 ;
        RECT 35.875 5.955 36.205 6.285 ;
        RECT 35.875 4.595 36.205 4.925 ;
        RECT 35.875 3.235 36.205 3.565 ;
        RECT 35.875 1.875 36.205 2.205 ;
        RECT 35.875 0.515 36.205 0.845 ;
        RECT 35.88 -8.32 36.2 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.235 15.475 37.565 15.805 ;
        RECT 37.235 10.035 37.565 10.365 ;
        RECT 37.235 8.675 37.565 9.005 ;
        RECT 37.235 7.315 37.565 7.645 ;
        RECT 37.235 5.955 37.565 6.285 ;
        RECT 37.235 4.595 37.565 4.925 ;
        RECT 37.235 3.235 37.565 3.565 ;
        RECT 37.235 1.875 37.565 2.205 ;
        RECT 37.235 0.515 37.565 0.845 ;
        RECT 37.24 -8.32 37.56 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.595 15.475 38.925 15.805 ;
        RECT 38.595 10.035 38.925 10.365 ;
        RECT 38.595 8.675 38.925 9.005 ;
        RECT 38.595 7.315 38.925 7.645 ;
        RECT 38.595 5.955 38.925 6.285 ;
        RECT 38.595 4.595 38.925 4.925 ;
        RECT 38.595 3.235 38.925 3.565 ;
        RECT 38.595 1.875 38.925 2.205 ;
        RECT 38.595 0.515 38.925 0.845 ;
        RECT 38.6 -8.32 38.92 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.955 15.475 40.285 15.805 ;
        RECT 39.955 11.395 40.285 11.725 ;
        RECT 39.955 10.035 40.285 10.365 ;
        RECT 39.955 8.675 40.285 9.005 ;
        RECT 39.955 7.315 40.285 7.645 ;
        RECT 39.955 5.955 40.285 6.285 ;
        RECT 39.955 4.595 40.285 4.925 ;
        RECT 39.955 3.235 40.285 3.565 ;
        RECT 39.955 1.875 40.285 2.205 ;
        RECT 39.955 0.515 40.285 0.845 ;
        RECT 39.96 -8.32 40.28 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.315 15.475 41.645 15.805 ;
        RECT 41.315 11.395 41.645 11.725 ;
        RECT 41.315 10.035 41.645 10.365 ;
        RECT 41.315 8.675 41.645 9.005 ;
        RECT 41.315 7.315 41.645 7.645 ;
        RECT 41.315 5.955 41.645 6.285 ;
        RECT 41.315 4.595 41.645 4.925 ;
        RECT 41.315 3.235 41.645 3.565 ;
        RECT 41.315 1.875 41.645 2.205 ;
        RECT 41.315 0.515 41.645 0.845 ;
        RECT 41.32 -8.32 41.64 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.675 15.475 43.005 15.805 ;
        RECT 42.675 11.395 43.005 11.725 ;
        RECT 42.675 10.035 43.005 10.365 ;
        RECT 42.675 8.675 43.005 9.005 ;
        RECT 42.675 7.315 43.005 7.645 ;
        RECT 42.675 5.955 43.005 6.285 ;
        RECT 42.675 4.595 43.005 4.925 ;
        RECT 42.675 3.235 43.005 3.565 ;
        RECT 42.675 1.875 43.005 2.205 ;
        RECT 42.675 0.515 43.005 0.845 ;
        RECT 42.68 -8.32 43 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.035 15.475 44.365 15.805 ;
        RECT 44.035 10.035 44.365 10.365 ;
        RECT 44.035 8.675 44.365 9.005 ;
        RECT 44.035 7.315 44.365 7.645 ;
        RECT 44.035 5.955 44.365 6.285 ;
        RECT 44.035 4.595 44.365 4.925 ;
        RECT 44.035 3.235 44.365 3.565 ;
        RECT 44.035 1.875 44.365 2.205 ;
        RECT 44.035 0.515 44.365 0.845 ;
        RECT 44.04 -8.32 44.36 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.395 15.475 45.725 15.805 ;
        RECT 45.395 10.035 45.725 10.365 ;
        RECT 45.395 8.675 45.725 9.005 ;
        RECT 45.395 7.315 45.725 7.645 ;
        RECT 45.395 5.955 45.725 6.285 ;
        RECT 45.395 4.595 45.725 4.925 ;
        RECT 45.395 3.235 45.725 3.565 ;
        RECT 45.395 1.875 45.725 2.205 ;
        RECT 45.395 0.515 45.725 0.845 ;
        RECT 45.4 -8.32 45.72 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.755 15.475 47.085 15.805 ;
        RECT 46.755 10.035 47.085 10.365 ;
        RECT 46.755 8.675 47.085 9.005 ;
        RECT 46.755 7.315 47.085 7.645 ;
        RECT 46.755 5.955 47.085 6.285 ;
        RECT 46.755 4.595 47.085 4.925 ;
        RECT 46.755 3.235 47.085 3.565 ;
        RECT 46.755 1.875 47.085 2.205 ;
        RECT 46.755 0.515 47.085 0.845 ;
        RECT 46.76 -8.32 47.08 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.115 15.475 48.445 15.805 ;
        RECT 48.115 10.035 48.445 10.365 ;
        RECT 48.115 8.675 48.445 9.005 ;
        RECT 48.115 7.315 48.445 7.645 ;
        RECT 48.115 5.955 48.445 6.285 ;
        RECT 48.115 4.595 48.445 4.925 ;
        RECT 48.115 3.235 48.445 3.565 ;
        RECT 48.115 1.875 48.445 2.205 ;
        RECT 48.115 0.515 48.445 0.845 ;
        RECT 48.12 -8.32 48.44 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.475 15.475 49.805 15.805 ;
        RECT 49.475 10.035 49.805 10.365 ;
        RECT 49.475 8.675 49.805 9.005 ;
        RECT 49.475 7.315 49.805 7.645 ;
        RECT 49.475 5.955 49.805 6.285 ;
        RECT 49.475 4.595 49.805 4.925 ;
        RECT 49.475 3.235 49.805 3.565 ;
        RECT 49.475 1.875 49.805 2.205 ;
        RECT 49.475 0.515 49.805 0.845 ;
        RECT 49.48 -8.32 49.8 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.835 15.475 51.165 15.805 ;
        RECT 50.835 11.395 51.165 11.725 ;
        RECT 50.835 10.035 51.165 10.365 ;
        RECT 50.835 8.675 51.165 9.005 ;
        RECT 50.835 7.315 51.165 7.645 ;
        RECT 50.835 5.955 51.165 6.285 ;
        RECT 50.835 4.595 51.165 4.925 ;
        RECT 50.835 3.235 51.165 3.565 ;
        RECT 50.835 1.875 51.165 2.205 ;
        RECT 50.835 0.515 51.165 0.845 ;
        RECT 50.84 -8.32 51.16 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.195 15.475 52.525 15.805 ;
        RECT 52.195 11.395 52.525 11.725 ;
        RECT 52.195 10.035 52.525 10.365 ;
        RECT 52.195 8.675 52.525 9.005 ;
        RECT 52.195 7.315 52.525 7.645 ;
        RECT 52.195 5.955 52.525 6.285 ;
        RECT 52.195 4.595 52.525 4.925 ;
        RECT 52.195 3.235 52.525 3.565 ;
        RECT 52.195 1.875 52.525 2.205 ;
        RECT 52.195 0.515 52.525 0.845 ;
        RECT 52.2 -8.32 52.52 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.555 15.475 53.885 15.805 ;
        RECT 53.555 11.395 53.885 11.725 ;
        RECT 53.555 10.035 53.885 10.365 ;
        RECT 53.555 8.675 53.885 9.005 ;
        RECT 53.555 7.315 53.885 7.645 ;
        RECT 53.555 5.955 53.885 6.285 ;
        RECT 53.555 4.595 53.885 4.925 ;
        RECT 53.555 3.235 53.885 3.565 ;
        RECT 53.555 1.875 53.885 2.205 ;
        RECT 53.555 0.515 53.885 0.845 ;
        RECT 53.56 -8.32 53.88 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.915 15.475 55.245 15.805 ;
        RECT 54.915 10.035 55.245 10.365 ;
        RECT 54.915 8.675 55.245 9.005 ;
        RECT 54.915 7.315 55.245 7.645 ;
        RECT 54.915 5.955 55.245 6.285 ;
        RECT 54.915 4.595 55.245 4.925 ;
        RECT 54.915 3.235 55.245 3.565 ;
        RECT 54.915 1.875 55.245 2.205 ;
        RECT 54.915 0.515 55.245 0.845 ;
        RECT 54.92 -8.32 55.24 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.275 15.475 56.605 15.805 ;
        RECT 56.275 10.035 56.605 10.365 ;
        RECT 56.275 8.675 56.605 9.005 ;
        RECT 56.275 7.315 56.605 7.645 ;
        RECT 56.275 5.955 56.605 6.285 ;
        RECT 56.275 4.595 56.605 4.925 ;
        RECT 56.275 3.235 56.605 3.565 ;
        RECT 56.275 1.875 56.605 2.205 ;
        RECT 56.275 0.515 56.605 0.845 ;
        RECT 56.28 -8.32 56.6 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.635 15.475 57.965 15.805 ;
        RECT 57.635 10.035 57.965 10.365 ;
        RECT 57.635 8.675 57.965 9.005 ;
        RECT 57.635 7.315 57.965 7.645 ;
        RECT 57.635 5.955 57.965 6.285 ;
        RECT 57.635 4.595 57.965 4.925 ;
        RECT 57.635 3.235 57.965 3.565 ;
        RECT 57.635 1.875 57.965 2.205 ;
        RECT 57.635 0.515 57.965 0.845 ;
        RECT 57.64 -8.32 57.96 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.995 15.475 59.325 15.805 ;
        RECT 58.995 10.035 59.325 10.365 ;
        RECT 58.995 8.675 59.325 9.005 ;
        RECT 58.995 7.315 59.325 7.645 ;
        RECT 58.995 5.955 59.325 6.285 ;
        RECT 58.995 4.595 59.325 4.925 ;
        RECT 58.995 3.235 59.325 3.565 ;
        RECT 58.995 1.875 59.325 2.205 ;
        RECT 58.995 0.515 59.325 0.845 ;
        RECT 59 -8.32 59.32 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.355 15.475 60.685 15.805 ;
        RECT 60.355 10.035 60.685 10.365 ;
        RECT 60.355 8.675 60.685 9.005 ;
        RECT 60.355 7.315 60.685 7.645 ;
        RECT 60.355 5.955 60.685 6.285 ;
        RECT 60.355 4.595 60.685 4.925 ;
        RECT 60.355 3.235 60.685 3.565 ;
        RECT 60.355 1.875 60.685 2.205 ;
        RECT 60.355 0.515 60.685 0.845 ;
        RECT 60.36 -8.32 60.68 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.715 15.475 62.045 15.805 ;
        RECT 61.715 10.035 62.045 10.365 ;
        RECT 61.715 8.675 62.045 9.005 ;
        RECT 61.715 7.315 62.045 7.645 ;
        RECT 61.715 5.955 62.045 6.285 ;
        RECT 61.715 4.595 62.045 4.925 ;
        RECT 61.715 3.235 62.045 3.565 ;
        RECT 61.715 1.875 62.045 2.205 ;
        RECT 61.715 0.515 62.045 0.845 ;
        RECT 61.72 -8.32 62.04 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.075 15.475 63.405 15.805 ;
        RECT 63.075 11.395 63.405 11.725 ;
        RECT 63.075 10.035 63.405 10.365 ;
        RECT 63.075 8.675 63.405 9.005 ;
        RECT 63.075 7.315 63.405 7.645 ;
        RECT 63.075 5.955 63.405 6.285 ;
        RECT 63.075 4.595 63.405 4.925 ;
        RECT 63.075 3.235 63.405 3.565 ;
        RECT 63.075 1.875 63.405 2.205 ;
        RECT 63.075 0.515 63.405 0.845 ;
        RECT 63.08 -8.32 63.4 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.435 15.475 64.765 15.805 ;
        RECT 64.435 11.395 64.765 11.725 ;
        RECT 64.435 10.035 64.765 10.365 ;
        RECT 64.435 8.675 64.765 9.005 ;
        RECT 64.435 7.315 64.765 7.645 ;
        RECT 64.435 5.955 64.765 6.285 ;
        RECT 64.435 4.595 64.765 4.925 ;
        RECT 64.435 3.235 64.765 3.565 ;
        RECT 64.435 1.875 64.765 2.205 ;
        RECT 64.435 0.515 64.765 0.845 ;
        RECT 64.44 -8.32 64.76 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.795 15.475 66.125 15.805 ;
        RECT 65.795 11.395 66.125 11.725 ;
        RECT 65.795 10.035 66.125 10.365 ;
        RECT 65.795 8.675 66.125 9.005 ;
        RECT 65.795 7.315 66.125 7.645 ;
        RECT 65.795 5.955 66.125 6.285 ;
        RECT 65.795 4.595 66.125 4.925 ;
        RECT 65.795 3.235 66.125 3.565 ;
        RECT 65.795 1.875 66.125 2.205 ;
        RECT 65.795 0.515 66.125 0.845 ;
        RECT 65.8 -8.32 66.12 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.155 15.475 67.485 15.805 ;
        RECT 67.155 10.035 67.485 10.365 ;
        RECT 67.155 8.675 67.485 9.005 ;
        RECT 67.155 7.315 67.485 7.645 ;
        RECT 67.155 5.955 67.485 6.285 ;
        RECT 67.155 4.595 67.485 4.925 ;
        RECT 67.155 3.235 67.485 3.565 ;
        RECT 67.155 1.875 67.485 2.205 ;
        RECT 67.155 0.515 67.485 0.845 ;
        RECT 67.16 -8.32 67.48 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.515 15.475 68.845 15.805 ;
        RECT 68.515 10.035 68.845 10.365 ;
        RECT 68.515 8.675 68.845 9.005 ;
        RECT 68.515 7.315 68.845 7.645 ;
        RECT 68.515 5.955 68.845 6.285 ;
        RECT 68.515 4.595 68.845 4.925 ;
        RECT 68.515 3.235 68.845 3.565 ;
        RECT 68.515 1.875 68.845 2.205 ;
        RECT 68.515 0.515 68.845 0.845 ;
        RECT 68.52 -8.32 68.84 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.875 15.475 70.205 15.805 ;
        RECT 69.875 10.035 70.205 10.365 ;
        RECT 69.875 8.675 70.205 9.005 ;
        RECT 69.875 7.315 70.205 7.645 ;
        RECT 69.875 5.955 70.205 6.285 ;
        RECT 69.875 4.595 70.205 4.925 ;
        RECT 69.875 3.235 70.205 3.565 ;
        RECT 69.875 1.875 70.205 2.205 ;
        RECT 69.875 0.515 70.205 0.845 ;
        RECT 69.88 -8.32 70.2 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.235 15.475 71.565 15.805 ;
        RECT 71.235 10.035 71.565 10.365 ;
        RECT 71.235 8.675 71.565 9.005 ;
        RECT 71.235 7.315 71.565 7.645 ;
        RECT 71.235 5.955 71.565 6.285 ;
        RECT 71.235 4.595 71.565 4.925 ;
        RECT 71.235 3.235 71.565 3.565 ;
        RECT 71.235 1.875 71.565 2.205 ;
        RECT 71.235 0.515 71.565 0.845 ;
        RECT 71.24 -8.32 71.56 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.595 15.475 72.925 15.805 ;
        RECT 72.595 10.035 72.925 10.365 ;
        RECT 72.595 8.675 72.925 9.005 ;
        RECT 72.595 7.315 72.925 7.645 ;
        RECT 72.595 5.955 72.925 6.285 ;
        RECT 72.595 4.595 72.925 4.925 ;
        RECT 72.595 3.235 72.925 3.565 ;
        RECT 72.595 1.875 72.925 2.205 ;
        RECT 72.595 0.515 72.925 0.845 ;
        RECT 72.6 -8.32 72.92 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 15.475 74.285 15.805 ;
        RECT 73.955 10.035 74.285 10.365 ;
        RECT 73.955 8.675 74.285 9.005 ;
        RECT 73.955 7.315 74.285 7.645 ;
        RECT 73.955 5.955 74.285 6.285 ;
        RECT 73.955 4.595 74.285 4.925 ;
        RECT 73.955 3.235 74.285 3.565 ;
        RECT 73.955 1.875 74.285 2.205 ;
        RECT 73.955 0.515 74.285 0.845 ;
        RECT 73.96 -8.32 74.28 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.315 15.475 75.645 15.805 ;
        RECT 75.315 11.395 75.645 11.725 ;
        RECT 75.315 10.035 75.645 10.365 ;
        RECT 75.315 8.675 75.645 9.005 ;
        RECT 75.315 7.315 75.645 7.645 ;
        RECT 75.315 5.955 75.645 6.285 ;
        RECT 75.315 4.595 75.645 4.925 ;
        RECT 75.315 3.235 75.645 3.565 ;
        RECT 75.315 1.875 75.645 2.205 ;
        RECT 75.315 0.515 75.645 0.845 ;
        RECT 75.32 -8.32 75.64 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 76.675 15.475 77.005 15.805 ;
        RECT 76.675 11.395 77.005 11.725 ;
        RECT 76.675 10.035 77.005 10.365 ;
        RECT 76.675 8.675 77.005 9.005 ;
        RECT 76.675 7.315 77.005 7.645 ;
        RECT 76.675 5.955 77.005 6.285 ;
        RECT 76.675 4.595 77.005 4.925 ;
        RECT 76.675 3.235 77.005 3.565 ;
        RECT 76.675 1.875 77.005 2.205 ;
        RECT 76.675 0.515 77.005 0.845 ;
        RECT 76.68 -8.32 77 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.035 15.475 78.365 15.805 ;
        RECT 78.035 11.395 78.365 11.725 ;
        RECT 78.035 10.035 78.365 10.365 ;
        RECT 78.035 8.675 78.365 9.005 ;
        RECT 78.035 7.315 78.365 7.645 ;
        RECT 78.035 5.955 78.365 6.285 ;
        RECT 78.035 4.595 78.365 4.925 ;
        RECT 78.035 3.235 78.365 3.565 ;
        RECT 78.035 1.875 78.365 2.205 ;
        RECT 78.035 0.515 78.365 0.845 ;
        RECT 78.04 -8.32 78.36 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 79.395 15.475 79.725 15.805 ;
        RECT 79.395 10.035 79.725 10.365 ;
        RECT 79.395 8.675 79.725 9.005 ;
        RECT 79.395 7.315 79.725 7.645 ;
        RECT 79.395 5.955 79.725 6.285 ;
        RECT 79.395 4.595 79.725 4.925 ;
        RECT 79.395 3.235 79.725 3.565 ;
        RECT 79.395 1.875 79.725 2.205 ;
        RECT 79.395 0.515 79.725 0.845 ;
        RECT 79.4 -8.32 79.72 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.755 15.475 81.085 15.805 ;
        RECT 80.755 10.035 81.085 10.365 ;
        RECT 80.755 8.675 81.085 9.005 ;
        RECT 80.755 7.315 81.085 7.645 ;
        RECT 80.755 5.955 81.085 6.285 ;
        RECT 80.755 4.595 81.085 4.925 ;
        RECT 80.755 3.235 81.085 3.565 ;
        RECT 80.755 1.875 81.085 2.205 ;
        RECT 80.755 0.515 81.085 0.845 ;
        RECT 80.76 -8.32 81.08 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.115 15.475 82.445 15.805 ;
        RECT 82.115 10.035 82.445 10.365 ;
        RECT 82.115 8.675 82.445 9.005 ;
        RECT 82.115 7.315 82.445 7.645 ;
        RECT 82.115 5.955 82.445 6.285 ;
        RECT 82.115 4.595 82.445 4.925 ;
        RECT 82.115 3.235 82.445 3.565 ;
        RECT 82.115 1.875 82.445 2.205 ;
        RECT 82.115 0.515 82.445 0.845 ;
        RECT 82.12 -8.32 82.44 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 83.475 15.475 83.805 15.805 ;
        RECT 83.475 10.035 83.805 10.365 ;
        RECT 83.475 8.675 83.805 9.005 ;
        RECT 83.475 7.315 83.805 7.645 ;
        RECT 83.475 5.955 83.805 6.285 ;
        RECT 83.475 4.595 83.805 4.925 ;
        RECT 83.475 3.235 83.805 3.565 ;
        RECT 83.475 1.875 83.805 2.205 ;
        RECT 83.475 0.515 83.805 0.845 ;
        RECT 83.48 -8.32 83.8 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.835 15.475 85.165 15.805 ;
        RECT 84.835 10.035 85.165 10.365 ;
        RECT 84.835 8.675 85.165 9.005 ;
        RECT 84.835 7.315 85.165 7.645 ;
        RECT 84.835 5.955 85.165 6.285 ;
        RECT 84.835 4.595 85.165 4.925 ;
        RECT 84.835 3.235 85.165 3.565 ;
        RECT 84.835 1.875 85.165 2.205 ;
        RECT 84.835 0.515 85.165 0.845 ;
        RECT 84.84 -8.32 85.16 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.195 15.475 86.525 15.805 ;
        RECT 86.195 10.035 86.525 10.365 ;
        RECT 86.195 8.675 86.525 9.005 ;
        RECT 86.195 7.315 86.525 7.645 ;
        RECT 86.195 5.955 86.525 6.285 ;
        RECT 86.195 4.595 86.525 4.925 ;
        RECT 86.195 3.235 86.525 3.565 ;
        RECT 86.195 1.875 86.525 2.205 ;
        RECT 86.195 0.515 86.525 0.845 ;
        RECT 86.2 -8.32 86.52 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.555 15.475 87.885 15.805 ;
        RECT 87.555 11.395 87.885 11.725 ;
        RECT 87.555 10.035 87.885 10.365 ;
        RECT 87.555 8.675 87.885 9.005 ;
        RECT 87.555 7.315 87.885 7.645 ;
        RECT 87.555 5.955 87.885 6.285 ;
        RECT 87.555 4.595 87.885 4.925 ;
        RECT 87.555 3.235 87.885 3.565 ;
        RECT 87.555 1.875 87.885 2.205 ;
        RECT 87.555 0.515 87.885 0.845 ;
        RECT 87.56 -8.32 87.88 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.915 15.475 89.245 15.805 ;
        RECT 88.915 11.395 89.245 11.725 ;
        RECT 88.915 10.035 89.245 10.365 ;
        RECT 88.915 8.675 89.245 9.005 ;
        RECT 88.915 7.315 89.245 7.645 ;
        RECT 88.915 5.955 89.245 6.285 ;
        RECT 88.915 4.595 89.245 4.925 ;
        RECT 88.915 3.235 89.245 3.565 ;
        RECT 88.915 1.875 89.245 2.205 ;
        RECT 88.915 0.515 89.245 0.845 ;
        RECT 88.92 -8.32 89.24 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.275 15.475 90.605 15.805 ;
        RECT 90.275 11.395 90.605 11.725 ;
        RECT 90.275 10.035 90.605 10.365 ;
        RECT 90.275 8.675 90.605 9.005 ;
        RECT 90.275 7.315 90.605 7.645 ;
        RECT 90.275 5.955 90.605 6.285 ;
        RECT 90.275 4.595 90.605 4.925 ;
        RECT 90.275 3.235 90.605 3.565 ;
        RECT 90.275 1.875 90.605 2.205 ;
        RECT 90.275 0.515 90.605 0.845 ;
        RECT 90.28 -8.32 90.6 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 91.635 15.475 91.965 15.805 ;
        RECT 91.635 10.035 91.965 10.365 ;
        RECT 91.635 8.675 91.965 9.005 ;
        RECT 91.635 7.315 91.965 7.645 ;
        RECT 91.635 5.955 91.965 6.285 ;
        RECT 91.635 4.595 91.965 4.925 ;
        RECT 91.635 3.235 91.965 3.565 ;
        RECT 91.635 1.875 91.965 2.205 ;
        RECT 91.635 0.515 91.965 0.845 ;
        RECT 91.64 -8.32 91.96 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.995 15.475 93.325 15.805 ;
        RECT 92.995 10.035 93.325 10.365 ;
        RECT 92.995 8.675 93.325 9.005 ;
        RECT 92.995 7.315 93.325 7.645 ;
        RECT 92.995 5.955 93.325 6.285 ;
        RECT 92.995 4.595 93.325 4.925 ;
        RECT 92.995 3.235 93.325 3.565 ;
        RECT 92.995 1.875 93.325 2.205 ;
        RECT 92.995 0.515 93.325 0.845 ;
        RECT 93 -8.32 93.32 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.355 15.475 94.685 15.805 ;
        RECT 94.355 10.035 94.685 10.365 ;
        RECT 94.355 8.675 94.685 9.005 ;
        RECT 94.355 7.315 94.685 7.645 ;
        RECT 94.355 5.955 94.685 6.285 ;
        RECT 94.355 4.595 94.685 4.925 ;
        RECT 94.355 3.235 94.685 3.565 ;
        RECT 94.355 1.875 94.685 2.205 ;
        RECT 94.355 0.515 94.685 0.845 ;
        RECT 94.36 -8.32 94.68 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.715 15.475 96.045 15.805 ;
        RECT 95.715 10.035 96.045 10.365 ;
        RECT 95.715 8.675 96.045 9.005 ;
        RECT 95.715 7.315 96.045 7.645 ;
        RECT 95.715 5.955 96.045 6.285 ;
        RECT 95.715 4.595 96.045 4.925 ;
        RECT 95.715 3.235 96.045 3.565 ;
        RECT 95.715 1.875 96.045 2.205 ;
        RECT 95.715 0.515 96.045 0.845 ;
        RECT 95.72 -8.32 96.04 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.075 15.475 97.405 15.805 ;
        RECT 97.075 10.035 97.405 10.365 ;
        RECT 97.075 8.675 97.405 9.005 ;
        RECT 97.075 7.315 97.405 7.645 ;
        RECT 97.075 5.955 97.405 6.285 ;
        RECT 97.075 4.595 97.405 4.925 ;
        RECT 97.075 3.235 97.405 3.565 ;
        RECT 97.075 1.875 97.405 2.205 ;
        RECT 97.075 0.515 97.405 0.845 ;
        RECT 97.08 -8.32 97.4 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.435 15.475 98.765 15.805 ;
        RECT 98.435 10.035 98.765 10.365 ;
        RECT 98.435 8.675 98.765 9.005 ;
        RECT 98.435 7.315 98.765 7.645 ;
        RECT 98.435 5.955 98.765 6.285 ;
        RECT 98.435 4.595 98.765 4.925 ;
        RECT 98.435 3.235 98.765 3.565 ;
        RECT 98.435 1.875 98.765 2.205 ;
        RECT 98.435 0.515 98.765 0.845 ;
        RECT 98.44 -8.32 98.76 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.795 15.475 100.125 15.805 ;
        RECT 99.795 11.395 100.125 11.725 ;
        RECT 99.795 10.035 100.125 10.365 ;
        RECT 99.795 8.675 100.125 9.005 ;
        RECT 99.795 7.315 100.125 7.645 ;
        RECT 99.795 5.955 100.125 6.285 ;
        RECT 99.795 4.595 100.125 4.925 ;
        RECT 99.795 3.235 100.125 3.565 ;
        RECT 99.795 1.875 100.125 2.205 ;
        RECT 99.795 0.515 100.125 0.845 ;
        RECT 99.8 -8.32 100.12 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.155 15.475 101.485 15.805 ;
        RECT 101.155 11.395 101.485 11.725 ;
        RECT 101.155 10.035 101.485 10.365 ;
        RECT 101.155 8.675 101.485 9.005 ;
        RECT 101.155 7.315 101.485 7.645 ;
        RECT 101.155 5.955 101.485 6.285 ;
        RECT 101.155 4.595 101.485 4.925 ;
        RECT 101.155 3.235 101.485 3.565 ;
        RECT 101.155 1.875 101.485 2.205 ;
        RECT 101.155 0.515 101.485 0.845 ;
        RECT 101.16 -8.32 101.48 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.515 15.475 102.845 15.805 ;
        RECT 102.515 11.395 102.845 11.725 ;
        RECT 102.515 10.035 102.845 10.365 ;
        RECT 102.515 8.675 102.845 9.005 ;
        RECT 102.515 7.315 102.845 7.645 ;
        RECT 102.515 5.955 102.845 6.285 ;
        RECT 102.515 4.595 102.845 4.925 ;
        RECT 102.515 3.235 102.845 3.565 ;
        RECT 102.515 1.875 102.845 2.205 ;
        RECT 102.515 0.515 102.845 0.845 ;
        RECT 102.52 -8.32 102.84 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.875 15.475 104.205 15.805 ;
        RECT 103.875 10.035 104.205 10.365 ;
        RECT 103.875 8.675 104.205 9.005 ;
        RECT 103.875 7.315 104.205 7.645 ;
        RECT 103.875 5.955 104.205 6.285 ;
        RECT 103.875 4.595 104.205 4.925 ;
        RECT 103.875 3.235 104.205 3.565 ;
        RECT 103.875 1.875 104.205 2.205 ;
        RECT 103.875 0.515 104.205 0.845 ;
        RECT 103.88 -8.32 104.2 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.235 15.475 105.565 15.805 ;
        RECT 105.235 10.035 105.565 10.365 ;
        RECT 105.235 8.675 105.565 9.005 ;
        RECT 105.235 7.315 105.565 7.645 ;
        RECT 105.235 5.955 105.565 6.285 ;
        RECT 105.235 4.595 105.565 4.925 ;
        RECT 105.235 3.235 105.565 3.565 ;
        RECT 105.235 1.875 105.565 2.205 ;
        RECT 105.235 0.515 105.565 0.845 ;
        RECT 105.24 -8.32 105.56 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.595 15.475 106.925 15.805 ;
        RECT 106.595 10.035 106.925 10.365 ;
        RECT 106.595 8.675 106.925 9.005 ;
        RECT 106.595 7.315 106.925 7.645 ;
        RECT 106.595 5.955 106.925 6.285 ;
        RECT 106.595 4.595 106.925 4.925 ;
        RECT 106.595 3.235 106.925 3.565 ;
        RECT 106.595 1.875 106.925 2.205 ;
        RECT 106.595 0.515 106.925 0.845 ;
        RECT 106.6 -8.32 106.92 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.955 15.475 108.285 15.805 ;
        RECT 107.955 10.035 108.285 10.365 ;
        RECT 107.955 8.675 108.285 9.005 ;
        RECT 107.955 7.315 108.285 7.645 ;
        RECT 107.955 5.955 108.285 6.285 ;
        RECT 107.955 4.595 108.285 4.925 ;
        RECT 107.955 3.235 108.285 3.565 ;
        RECT 107.955 1.875 108.285 2.205 ;
        RECT 107.955 0.515 108.285 0.845 ;
        RECT 107.96 -8.32 108.28 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.315 15.475 109.645 15.805 ;
        RECT 109.315 10.035 109.645 10.365 ;
        RECT 109.315 8.675 109.645 9.005 ;
        RECT 109.315 7.315 109.645 7.645 ;
        RECT 109.315 5.955 109.645 6.285 ;
        RECT 109.315 4.595 109.645 4.925 ;
        RECT 109.315 3.235 109.645 3.565 ;
        RECT 109.315 1.875 109.645 2.205 ;
        RECT 109.315 0.515 109.645 0.845 ;
        RECT 109.32 -8.32 109.64 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.675 15.475 111.005 15.805 ;
        RECT 110.675 10.035 111.005 10.365 ;
        RECT 110.675 8.675 111.005 9.005 ;
        RECT 110.675 7.315 111.005 7.645 ;
        RECT 110.675 5.955 111.005 6.285 ;
        RECT 110.675 4.595 111.005 4.925 ;
        RECT 110.675 3.235 111.005 3.565 ;
        RECT 110.675 1.875 111.005 2.205 ;
        RECT 110.675 0.515 111.005 0.845 ;
        RECT 110.68 -8.32 111 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.035 15.475 112.365 15.805 ;
        RECT 112.035 11.395 112.365 11.725 ;
        RECT 112.035 10.035 112.365 10.365 ;
        RECT 112.035 8.675 112.365 9.005 ;
        RECT 112.035 7.315 112.365 7.645 ;
        RECT 112.035 5.955 112.365 6.285 ;
        RECT 112.035 4.595 112.365 4.925 ;
        RECT 112.035 3.235 112.365 3.565 ;
        RECT 112.035 1.875 112.365 2.205 ;
        RECT 112.035 0.515 112.365 0.845 ;
        RECT 112.04 -8.32 112.36 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.395 4.595 113.725 4.925 ;
        RECT 113.395 3.235 113.725 3.565 ;
        RECT 113.395 1.875 113.725 2.205 ;
        RECT 113.395 0.515 113.725 0.845 ;
        RECT 113.4 -8.32 113.72 15.805 ;
        RECT 113.395 15.475 113.725 15.805 ;
        RECT 113.395 11.395 113.725 11.725 ;
        RECT 113.395 10.035 113.725 10.365 ;
        RECT 113.395 8.675 113.725 9.005 ;
        RECT 113.395 7.315 113.725 7.645 ;
        RECT 113.395 5.955 113.725 6.285 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 634.955 10.715 635.285 11.045 ;
        RECT 634.955 9.355 635.285 9.685 ;
        RECT 634.955 7.995 635.285 8.325 ;
        RECT 634.955 6.635 635.285 6.965 ;
        RECT 634.955 5.275 635.285 5.605 ;
        RECT 634.955 3.915 635.285 4.245 ;
        RECT 634.955 2.555 635.285 2.885 ;
        RECT 634.955 1.195 635.285 1.525 ;
        RECT 634.955 -0.165 635.285 0.165 ;
        RECT 634.96 -8.32 635.28 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 636.315 10.715 636.645 11.045 ;
        RECT 636.315 9.355 636.645 9.685 ;
        RECT 636.315 7.995 636.645 8.325 ;
        RECT 636.315 6.635 636.645 6.965 ;
        RECT 636.315 5.275 636.645 5.605 ;
        RECT 636.315 3.915 636.645 4.245 ;
        RECT 636.315 2.555 636.645 2.885 ;
        RECT 636.315 1.195 636.645 1.525 ;
        RECT 636.315 -0.165 636.645 0.165 ;
        RECT 636.32 -8.32 636.64 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 637.675 10.715 638.005 11.045 ;
        RECT 637.675 9.355 638.005 9.685 ;
        RECT 637.675 7.995 638.005 8.325 ;
        RECT 637.675 6.635 638.005 6.965 ;
        RECT 637.675 5.275 638.005 5.605 ;
        RECT 637.675 3.915 638.005 4.245 ;
        RECT 637.675 2.555 638.005 2.885 ;
        RECT 637.675 1.195 638.005 1.525 ;
        RECT 637.675 -0.165 638.005 0.165 ;
        RECT 637.68 -8.32 638 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 639.035 10.715 639.365 11.045 ;
        RECT 639.035 9.355 639.365 9.685 ;
        RECT 639.035 7.995 639.365 8.325 ;
        RECT 639.035 6.635 639.365 6.965 ;
        RECT 639.035 5.275 639.365 5.605 ;
        RECT 639.035 3.915 639.365 4.245 ;
        RECT 639.035 2.555 639.365 2.885 ;
        RECT 639.035 1.195 639.365 1.525 ;
        RECT 639.035 -0.165 639.365 0.165 ;
        RECT 639.04 -8.32 639.36 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 640.395 10.715 640.725 11.045 ;
        RECT 640.395 9.355 640.725 9.685 ;
        RECT 640.395 7.995 640.725 8.325 ;
        RECT 640.395 6.635 640.725 6.965 ;
        RECT 640.395 5.275 640.725 5.605 ;
        RECT 640.395 3.915 640.725 4.245 ;
        RECT 640.395 2.555 640.725 2.885 ;
        RECT 640.395 1.195 640.725 1.525 ;
        RECT 640.395 -0.165 640.725 0.165 ;
        RECT 640.4 -8.32 640.72 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 641.755 10.715 642.085 11.045 ;
        RECT 641.755 9.355 642.085 9.685 ;
        RECT 641.755 7.995 642.085 8.325 ;
        RECT 641.755 6.635 642.085 6.965 ;
        RECT 641.755 5.275 642.085 5.605 ;
        RECT 641.755 3.915 642.085 4.245 ;
        RECT 641.755 2.555 642.085 2.885 ;
        RECT 641.755 1.195 642.085 1.525 ;
        RECT 641.755 -0.165 642.085 0.165 ;
        RECT 641.76 -8.32 642.08 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 643.115 10.715 643.445 11.045 ;
        RECT 643.115 9.355 643.445 9.685 ;
        RECT 643.115 7.995 643.445 8.325 ;
        RECT 643.115 6.635 643.445 6.965 ;
        RECT 643.115 5.275 643.445 5.605 ;
        RECT 643.115 3.915 643.445 4.245 ;
        RECT 643.115 2.555 643.445 2.885 ;
        RECT 643.115 1.195 643.445 1.525 ;
        RECT 643.115 -0.165 643.445 0.165 ;
        RECT 643.12 -8.32 643.44 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 644.475 10.715 644.805 11.045 ;
        RECT 644.475 9.355 644.805 9.685 ;
        RECT 644.475 7.995 644.805 8.325 ;
        RECT 644.475 6.635 644.805 6.965 ;
        RECT 644.475 5.275 644.805 5.605 ;
        RECT 644.475 3.915 644.805 4.245 ;
        RECT 644.475 2.555 644.805 2.885 ;
        RECT 644.475 1.195 644.805 1.525 ;
        RECT 644.475 -0.165 644.805 0.165 ;
        RECT 644.48 -8.32 644.8 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 645.835 10.715 646.165 11.045 ;
        RECT 645.835 9.355 646.165 9.685 ;
        RECT 645.835 7.995 646.165 8.325 ;
        RECT 645.835 6.635 646.165 6.965 ;
        RECT 645.835 5.275 646.165 5.605 ;
        RECT 645.835 3.915 646.165 4.245 ;
        RECT 645.835 2.555 646.165 2.885 ;
        RECT 645.835 1.195 646.165 1.525 ;
        RECT 645.835 -0.165 646.165 0.165 ;
        RECT 645.84 -8.32 646.16 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 647.195 10.715 647.525 11.045 ;
        RECT 647.195 9.355 647.525 9.685 ;
        RECT 647.195 7.995 647.525 8.325 ;
        RECT 647.195 6.635 647.525 6.965 ;
        RECT 647.195 5.275 647.525 5.605 ;
        RECT 647.195 3.915 647.525 4.245 ;
        RECT 647.195 2.555 647.525 2.885 ;
        RECT 647.195 1.195 647.525 1.525 ;
        RECT 647.195 -0.165 647.525 0.165 ;
        RECT 647.2 -8.32 647.52 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 648.555 10.715 648.885 11.045 ;
        RECT 648.555 9.355 648.885 9.685 ;
        RECT 648.555 7.995 648.885 8.325 ;
        RECT 648.555 6.635 648.885 6.965 ;
        RECT 648.555 5.275 648.885 5.605 ;
        RECT 648.555 3.915 648.885 4.245 ;
        RECT 648.555 2.555 648.885 2.885 ;
        RECT 648.555 1.195 648.885 1.525 ;
        RECT 648.555 -0.165 648.885 0.165 ;
        RECT 648.56 -8.32 648.88 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 649.915 10.715 650.245 11.045 ;
        RECT 649.915 9.355 650.245 9.685 ;
        RECT 649.915 7.995 650.245 8.325 ;
        RECT 649.915 6.635 650.245 6.965 ;
        RECT 649.915 5.275 650.245 5.605 ;
        RECT 649.915 3.915 650.245 4.245 ;
        RECT 649.915 2.555 650.245 2.885 ;
        RECT 649.915 1.195 650.245 1.525 ;
        RECT 649.915 -0.165 650.245 0.165 ;
        RECT 649.92 -8.32 650.24 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 651.275 10.715 651.605 11.045 ;
        RECT 651.275 9.355 651.605 9.685 ;
        RECT 651.275 7.995 651.605 8.325 ;
        RECT 651.275 6.635 651.605 6.965 ;
        RECT 651.275 5.275 651.605 5.605 ;
        RECT 651.275 3.915 651.605 4.245 ;
        RECT 651.275 2.555 651.605 2.885 ;
        RECT 651.275 1.195 651.605 1.525 ;
        RECT 651.275 -0.165 651.605 0.165 ;
        RECT 651.28 -8.32 651.6 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 652.635 10.715 652.965 11.045 ;
        RECT 652.635 9.355 652.965 9.685 ;
        RECT 652.635 7.995 652.965 8.325 ;
        RECT 652.635 6.635 652.965 6.965 ;
        RECT 652.635 5.275 652.965 5.605 ;
        RECT 652.635 3.915 652.965 4.245 ;
        RECT 652.635 2.555 652.965 2.885 ;
        RECT 652.635 1.195 652.965 1.525 ;
        RECT 652.635 -0.165 652.965 0.165 ;
        RECT 652.64 -8.32 652.96 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 653.995 10.715 654.325 11.045 ;
        RECT 653.995 9.355 654.325 9.685 ;
        RECT 653.995 7.995 654.325 8.325 ;
        RECT 653.995 6.635 654.325 6.965 ;
        RECT 653.995 5.275 654.325 5.605 ;
        RECT 653.995 3.915 654.325 4.245 ;
        RECT 653.995 2.555 654.325 2.885 ;
        RECT 653.995 1.195 654.325 1.525 ;
        RECT 653.995 -0.165 654.325 0.165 ;
        RECT 654 -8.32 654.32 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 655.355 10.715 655.685 11.045 ;
        RECT 655.355 9.355 655.685 9.685 ;
        RECT 655.355 7.995 655.685 8.325 ;
        RECT 655.355 6.635 655.685 6.965 ;
        RECT 655.355 5.275 655.685 5.605 ;
        RECT 655.355 3.915 655.685 4.245 ;
        RECT 655.355 2.555 655.685 2.885 ;
        RECT 655.355 1.195 655.685 1.525 ;
        RECT 655.355 -0.165 655.685 0.165 ;
        RECT 655.36 -8.32 655.68 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 656.715 10.715 657.045 11.045 ;
        RECT 656.715 9.355 657.045 9.685 ;
        RECT 656.715 7.995 657.045 8.325 ;
        RECT 656.715 6.635 657.045 6.965 ;
        RECT 656.715 5.275 657.045 5.605 ;
        RECT 656.715 3.915 657.045 4.245 ;
        RECT 656.715 2.555 657.045 2.885 ;
        RECT 656.715 1.195 657.045 1.525 ;
        RECT 656.715 -0.165 657.045 0.165 ;
        RECT 656.72 -8.32 657.04 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 658.075 10.715 658.405 11.045 ;
        RECT 658.075 9.355 658.405 9.685 ;
        RECT 658.075 7.995 658.405 8.325 ;
        RECT 658.075 6.635 658.405 6.965 ;
        RECT 658.075 5.275 658.405 5.605 ;
        RECT 658.075 3.915 658.405 4.245 ;
        RECT 658.075 2.555 658.405 2.885 ;
        RECT 658.075 1.195 658.405 1.525 ;
        RECT 658.075 -0.165 658.405 0.165 ;
        RECT 658.08 -8.32 658.4 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 659.435 10.715 659.765 11.045 ;
        RECT 659.435 9.355 659.765 9.685 ;
        RECT 659.435 7.995 659.765 8.325 ;
        RECT 659.435 6.635 659.765 6.965 ;
        RECT 659.435 5.275 659.765 5.605 ;
        RECT 659.435 3.915 659.765 4.245 ;
        RECT 659.435 2.555 659.765 2.885 ;
        RECT 659.435 1.195 659.765 1.525 ;
        RECT 659.435 -0.165 659.765 0.165 ;
        RECT 659.44 -8.32 659.76 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 660.795 10.715 661.125 11.045 ;
        RECT 660.795 9.355 661.125 9.685 ;
        RECT 660.795 7.995 661.125 8.325 ;
        RECT 660.795 6.635 661.125 6.965 ;
        RECT 660.795 5.275 661.125 5.605 ;
        RECT 660.795 3.915 661.125 4.245 ;
        RECT 660.795 2.555 661.125 2.885 ;
        RECT 660.795 1.195 661.125 1.525 ;
        RECT 660.795 -0.165 661.125 0.165 ;
        RECT 660.8 -8.32 661.12 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 662.155 10.715 662.485 11.045 ;
        RECT 662.155 9.355 662.485 9.685 ;
        RECT 662.155 7.995 662.485 8.325 ;
        RECT 662.155 6.635 662.485 6.965 ;
        RECT 662.155 5.275 662.485 5.605 ;
        RECT 662.155 3.915 662.485 4.245 ;
        RECT 662.155 2.555 662.485 2.885 ;
        RECT 662.155 1.195 662.485 1.525 ;
        RECT 662.155 -0.165 662.485 0.165 ;
        RECT 662.16 -8.32 662.48 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 663.515 10.715 663.845 11.045 ;
        RECT 663.515 9.355 663.845 9.685 ;
        RECT 663.515 7.995 663.845 8.325 ;
        RECT 663.515 6.635 663.845 6.965 ;
        RECT 663.515 5.275 663.845 5.605 ;
        RECT 663.515 3.915 663.845 4.245 ;
        RECT 663.515 2.555 663.845 2.885 ;
        RECT 663.515 1.195 663.845 1.525 ;
        RECT 663.515 -0.165 663.845 0.165 ;
        RECT 663.52 -8.32 663.84 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 664.875 10.715 665.205 11.045 ;
        RECT 664.875 9.355 665.205 9.685 ;
        RECT 664.875 7.995 665.205 8.325 ;
        RECT 664.875 6.635 665.205 6.965 ;
        RECT 664.875 5.275 665.205 5.605 ;
        RECT 664.875 3.915 665.205 4.245 ;
        RECT 664.875 2.555 665.205 2.885 ;
        RECT 664.875 1.195 665.205 1.525 ;
        RECT 664.875 -0.165 665.205 0.165 ;
        RECT 664.88 -8.32 665.2 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 666.235 10.715 666.565 11.045 ;
        RECT 666.235 9.355 666.565 9.685 ;
        RECT 666.235 7.995 666.565 8.325 ;
        RECT 666.235 6.635 666.565 6.965 ;
        RECT 666.235 5.275 666.565 5.605 ;
        RECT 666.235 3.915 666.565 4.245 ;
        RECT 666.235 2.555 666.565 2.885 ;
        RECT 666.235 1.195 666.565 1.525 ;
        RECT 666.235 -0.165 666.565 0.165 ;
        RECT 666.24 -8.32 666.56 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 667.595 10.715 667.925 11.045 ;
        RECT 667.595 9.355 667.925 9.685 ;
        RECT 667.595 7.995 667.925 8.325 ;
        RECT 667.595 6.635 667.925 6.965 ;
        RECT 667.595 5.275 667.925 5.605 ;
        RECT 667.595 3.915 667.925 4.245 ;
        RECT 667.595 2.555 667.925 2.885 ;
        RECT 667.595 1.195 667.925 1.525 ;
        RECT 667.595 -0.165 667.925 0.165 ;
        RECT 667.6 -8.32 667.92 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 668.955 10.715 669.285 11.045 ;
        RECT 668.955 9.355 669.285 9.685 ;
        RECT 668.955 7.995 669.285 8.325 ;
        RECT 668.955 6.635 669.285 6.965 ;
        RECT 668.955 5.275 669.285 5.605 ;
        RECT 668.955 3.915 669.285 4.245 ;
        RECT 668.955 2.555 669.285 2.885 ;
        RECT 668.955 1.195 669.285 1.525 ;
        RECT 668.955 -0.165 669.285 0.165 ;
        RECT 668.96 -8.32 669.28 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 670.315 10.715 670.645 11.045 ;
        RECT 670.315 9.355 670.645 9.685 ;
        RECT 670.315 7.995 670.645 8.325 ;
        RECT 670.315 6.635 670.645 6.965 ;
        RECT 670.315 5.275 670.645 5.605 ;
        RECT 670.315 3.915 670.645 4.245 ;
        RECT 670.315 2.555 670.645 2.885 ;
        RECT 670.315 1.195 670.645 1.525 ;
        RECT 670.315 -0.165 670.645 0.165 ;
        RECT 670.32 -8.32 670.64 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 671.675 10.715 672.005 11.045 ;
        RECT 671.675 9.355 672.005 9.685 ;
        RECT 671.675 7.995 672.005 8.325 ;
        RECT 671.675 6.635 672.005 6.965 ;
        RECT 671.675 5.275 672.005 5.605 ;
        RECT 671.675 3.915 672.005 4.245 ;
        RECT 671.675 2.555 672.005 2.885 ;
        RECT 671.675 1.195 672.005 1.525 ;
        RECT 671.675 -0.165 672.005 0.165 ;
        RECT 671.68 -8.32 672 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 673.035 10.715 673.365 11.045 ;
        RECT 673.035 9.355 673.365 9.685 ;
        RECT 673.035 7.995 673.365 8.325 ;
        RECT 673.035 6.635 673.365 6.965 ;
        RECT 673.035 5.275 673.365 5.605 ;
        RECT 673.035 3.915 673.365 4.245 ;
        RECT 673.035 2.555 673.365 2.885 ;
        RECT 673.035 1.195 673.365 1.525 ;
        RECT 673.035 -0.165 673.365 0.165 ;
        RECT 673.04 -8.32 673.36 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 674.395 10.715 674.725 11.045 ;
        RECT 674.395 9.355 674.725 9.685 ;
        RECT 674.395 7.995 674.725 8.325 ;
        RECT 674.395 6.635 674.725 6.965 ;
        RECT 674.395 5.275 674.725 5.605 ;
        RECT 674.395 3.915 674.725 4.245 ;
        RECT 674.395 2.555 674.725 2.885 ;
        RECT 674.395 1.195 674.725 1.525 ;
        RECT 674.395 -0.165 674.725 0.165 ;
        RECT 674.4 -8.32 674.72 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 675.755 10.715 676.085 11.045 ;
        RECT 675.755 9.355 676.085 9.685 ;
        RECT 675.755 7.995 676.085 8.325 ;
        RECT 675.755 6.635 676.085 6.965 ;
        RECT 675.755 5.275 676.085 5.605 ;
        RECT 675.755 3.915 676.085 4.245 ;
        RECT 675.755 2.555 676.085 2.885 ;
        RECT 675.755 1.195 676.085 1.525 ;
        RECT 675.755 -0.165 676.085 0.165 ;
        RECT 675.76 -8.32 676.08 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 677.115 10.715 677.445 11.045 ;
        RECT 677.115 9.355 677.445 9.685 ;
        RECT 677.115 7.995 677.445 8.325 ;
        RECT 677.115 6.635 677.445 6.965 ;
        RECT 677.115 5.275 677.445 5.605 ;
        RECT 677.115 3.915 677.445 4.245 ;
        RECT 677.115 2.555 677.445 2.885 ;
        RECT 677.115 1.195 677.445 1.525 ;
        RECT 677.115 -0.165 677.445 0.165 ;
        RECT 677.12 -8.32 677.44 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 678.475 10.715 678.805 11.045 ;
        RECT 678.475 9.355 678.805 9.685 ;
        RECT 678.475 7.995 678.805 8.325 ;
        RECT 678.475 6.635 678.805 6.965 ;
        RECT 678.475 5.275 678.805 5.605 ;
        RECT 678.475 3.915 678.805 4.245 ;
        RECT 678.475 2.555 678.805 2.885 ;
        RECT 678.475 1.195 678.805 1.525 ;
        RECT 678.475 -0.165 678.805 0.165 ;
        RECT 678.48 -8.32 678.8 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 679.835 10.715 680.165 11.045 ;
        RECT 679.835 9.355 680.165 9.685 ;
        RECT 679.835 7.995 680.165 8.325 ;
        RECT 679.835 6.635 680.165 6.965 ;
        RECT 679.835 5.275 680.165 5.605 ;
        RECT 679.835 3.915 680.165 4.245 ;
        RECT 679.835 2.555 680.165 2.885 ;
        RECT 679.835 1.195 680.165 1.525 ;
        RECT 679.835 -0.165 680.165 0.165 ;
        RECT 679.84 -8.32 680.16 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 681.195 10.715 681.525 11.045 ;
        RECT 681.195 9.355 681.525 9.685 ;
        RECT 681.195 7.995 681.525 8.325 ;
        RECT 681.195 6.635 681.525 6.965 ;
        RECT 681.195 5.275 681.525 5.605 ;
        RECT 681.195 3.915 681.525 4.245 ;
        RECT 681.195 2.555 681.525 2.885 ;
        RECT 681.195 1.195 681.525 1.525 ;
        RECT 681.195 -0.165 681.525 0.165 ;
        RECT 681.2 -8.32 681.52 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 682.555 10.715 682.885 11.045 ;
        RECT 682.555 9.355 682.885 9.685 ;
        RECT 682.555 7.995 682.885 8.325 ;
        RECT 682.555 6.635 682.885 6.965 ;
        RECT 682.555 5.275 682.885 5.605 ;
        RECT 682.555 3.915 682.885 4.245 ;
        RECT 682.555 2.555 682.885 2.885 ;
        RECT 682.555 1.195 682.885 1.525 ;
        RECT 682.555 -0.165 682.885 0.165 ;
        RECT 682.56 -8.32 682.88 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 683.915 10.715 684.245 11.045 ;
        RECT 683.915 9.355 684.245 9.685 ;
        RECT 683.915 7.995 684.245 8.325 ;
        RECT 683.915 6.635 684.245 6.965 ;
        RECT 683.915 5.275 684.245 5.605 ;
        RECT 683.915 3.915 684.245 4.245 ;
        RECT 683.915 2.555 684.245 2.885 ;
        RECT 683.915 1.195 684.245 1.525 ;
        RECT 683.915 -0.165 684.245 0.165 ;
        RECT 683.92 -8.32 684.24 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 685.275 10.715 685.605 11.045 ;
        RECT 685.275 9.355 685.605 9.685 ;
        RECT 685.275 7.995 685.605 8.325 ;
        RECT 685.275 6.635 685.605 6.965 ;
        RECT 685.275 5.275 685.605 5.605 ;
        RECT 685.275 3.915 685.605 4.245 ;
        RECT 685.275 2.555 685.605 2.885 ;
        RECT 685.275 1.195 685.605 1.525 ;
        RECT 685.275 -0.165 685.605 0.165 ;
        RECT 685.28 -8.32 685.6 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 686.635 10.715 686.965 11.045 ;
        RECT 686.635 9.355 686.965 9.685 ;
        RECT 686.635 7.995 686.965 8.325 ;
        RECT 686.635 6.635 686.965 6.965 ;
        RECT 686.635 5.275 686.965 5.605 ;
        RECT 686.635 3.915 686.965 4.245 ;
        RECT 686.635 2.555 686.965 2.885 ;
        RECT 686.635 1.195 686.965 1.525 ;
        RECT 686.635 -0.165 686.965 0.165 ;
        RECT 686.64 -8.32 686.96 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 687.995 10.715 688.325 11.045 ;
        RECT 687.995 9.355 688.325 9.685 ;
        RECT 687.995 7.995 688.325 8.325 ;
        RECT 687.995 6.635 688.325 6.965 ;
        RECT 687.995 5.275 688.325 5.605 ;
        RECT 687.995 3.915 688.325 4.245 ;
        RECT 687.995 2.555 688.325 2.885 ;
        RECT 687.995 1.195 688.325 1.525 ;
        RECT 687.995 -0.165 688.325 0.165 ;
        RECT 688 -8.32 688.32 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 689.355 10.715 689.685 11.045 ;
        RECT 689.355 9.355 689.685 9.685 ;
        RECT 689.355 7.995 689.685 8.325 ;
        RECT 689.355 6.635 689.685 6.965 ;
        RECT 689.355 5.275 689.685 5.605 ;
        RECT 689.355 3.915 689.685 4.245 ;
        RECT 689.355 2.555 689.685 2.885 ;
        RECT 689.355 1.195 689.685 1.525 ;
        RECT 689.355 -0.165 689.685 0.165 ;
        RECT 689.36 -8.32 689.68 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 690.715 10.715 691.045 11.045 ;
        RECT 690.715 9.355 691.045 9.685 ;
        RECT 690.715 7.995 691.045 8.325 ;
        RECT 690.715 6.635 691.045 6.965 ;
        RECT 690.715 5.275 691.045 5.605 ;
        RECT 690.715 3.915 691.045 4.245 ;
        RECT 690.715 2.555 691.045 2.885 ;
        RECT 690.715 1.195 691.045 1.525 ;
        RECT 690.715 -0.165 691.045 0.165 ;
        RECT 690.72 -8.32 691.04 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 692.075 10.715 692.405 11.045 ;
        RECT 692.075 9.355 692.405 9.685 ;
        RECT 692.075 7.995 692.405 8.325 ;
        RECT 692.075 6.635 692.405 6.965 ;
        RECT 692.075 5.275 692.405 5.605 ;
        RECT 692.075 3.915 692.405 4.245 ;
        RECT 692.075 2.555 692.405 2.885 ;
        RECT 692.075 1.195 692.405 1.525 ;
        RECT 692.075 -0.165 692.405 0.165 ;
        RECT 692.08 -8.32 692.4 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 693.435 10.715 693.765 11.045 ;
        RECT 693.435 9.355 693.765 9.685 ;
        RECT 693.435 7.995 693.765 8.325 ;
        RECT 693.435 6.635 693.765 6.965 ;
        RECT 693.435 5.275 693.765 5.605 ;
        RECT 693.435 3.915 693.765 4.245 ;
        RECT 693.435 2.555 693.765 2.885 ;
        RECT 693.435 1.195 693.765 1.525 ;
        RECT 693.435 -0.165 693.765 0.165 ;
        RECT 693.44 -8.32 693.76 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 694.795 10.715 695.125 11.045 ;
        RECT 694.795 9.355 695.125 9.685 ;
        RECT 694.795 7.995 695.125 8.325 ;
        RECT 694.795 6.635 695.125 6.965 ;
        RECT 694.795 5.275 695.125 5.605 ;
        RECT 694.795 3.915 695.125 4.245 ;
        RECT 694.795 2.555 695.125 2.885 ;
        RECT 694.795 1.195 695.125 1.525 ;
        RECT 694.795 -0.165 695.125 0.165 ;
        RECT 694.8 -8.32 695.12 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 696.155 10.715 696.485 11.045 ;
        RECT 696.155 9.355 696.485 9.685 ;
        RECT 696.155 7.995 696.485 8.325 ;
        RECT 696.155 6.635 696.485 6.965 ;
        RECT 696.155 5.275 696.485 5.605 ;
        RECT 696.155 3.915 696.485 4.245 ;
        RECT 696.155 2.555 696.485 2.885 ;
        RECT 696.155 1.195 696.485 1.525 ;
        RECT 696.155 -0.165 696.485 0.165 ;
        RECT 696.16 -8.32 696.48 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 697.515 10.715 697.845 11.045 ;
        RECT 697.515 9.355 697.845 9.685 ;
        RECT 697.515 7.995 697.845 8.325 ;
        RECT 697.515 6.635 697.845 6.965 ;
        RECT 697.515 5.275 697.845 5.605 ;
        RECT 697.515 3.915 697.845 4.245 ;
        RECT 697.515 2.555 697.845 2.885 ;
        RECT 697.515 1.195 697.845 1.525 ;
        RECT 697.515 -0.165 697.845 0.165 ;
        RECT 697.52 -8.32 697.84 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 698.875 10.715 699.205 11.045 ;
        RECT 698.875 9.355 699.205 9.685 ;
        RECT 698.875 7.995 699.205 8.325 ;
        RECT 698.875 6.635 699.205 6.965 ;
        RECT 698.875 5.275 699.205 5.605 ;
        RECT 698.875 3.915 699.205 4.245 ;
        RECT 698.875 2.555 699.205 2.885 ;
        RECT 698.875 1.195 699.205 1.525 ;
        RECT 698.875 -0.165 699.205 0.165 ;
        RECT 698.88 -8.32 699.2 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 700.235 10.715 700.565 11.045 ;
        RECT 700.235 9.355 700.565 9.685 ;
        RECT 700.235 7.995 700.565 8.325 ;
        RECT 700.235 6.635 700.565 6.965 ;
        RECT 700.235 5.275 700.565 5.605 ;
        RECT 700.235 3.915 700.565 4.245 ;
        RECT 700.235 2.555 700.565 2.885 ;
        RECT 700.235 1.195 700.565 1.525 ;
        RECT 700.235 -0.165 700.565 0.165 ;
        RECT 700.24 -8.32 700.56 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 701.595 10.715 701.925 11.045 ;
        RECT 701.595 9.355 701.925 9.685 ;
        RECT 701.595 7.995 701.925 8.325 ;
        RECT 701.595 6.635 701.925 6.965 ;
        RECT 701.595 5.275 701.925 5.605 ;
        RECT 701.595 3.915 701.925 4.245 ;
        RECT 701.595 2.555 701.925 2.885 ;
        RECT 701.595 1.195 701.925 1.525 ;
        RECT 701.595 -0.165 701.925 0.165 ;
        RECT 701.6 -8.32 701.92 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 702.955 10.715 703.285 11.045 ;
        RECT 702.955 9.355 703.285 9.685 ;
        RECT 702.955 7.995 703.285 8.325 ;
        RECT 702.955 6.635 703.285 6.965 ;
        RECT 702.955 5.275 703.285 5.605 ;
        RECT 702.955 3.915 703.285 4.245 ;
        RECT 702.955 2.555 703.285 2.885 ;
        RECT 702.955 1.195 703.285 1.525 ;
        RECT 702.955 -0.165 703.285 0.165 ;
        RECT 702.96 -8.32 703.28 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 704.315 10.715 704.645 11.045 ;
        RECT 704.315 9.355 704.645 9.685 ;
        RECT 704.315 7.995 704.645 8.325 ;
        RECT 704.315 6.635 704.645 6.965 ;
        RECT 704.315 5.275 704.645 5.605 ;
        RECT 704.315 3.915 704.645 4.245 ;
        RECT 704.315 2.555 704.645 2.885 ;
        RECT 704.315 1.195 704.645 1.525 ;
        RECT 704.315 -0.165 704.645 0.165 ;
        RECT 704.32 -8.32 704.64 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 705.675 10.715 706.005 11.045 ;
        RECT 705.675 9.355 706.005 9.685 ;
        RECT 705.675 7.995 706.005 8.325 ;
        RECT 705.675 6.635 706.005 6.965 ;
        RECT 705.675 5.275 706.005 5.605 ;
        RECT 705.675 3.915 706.005 4.245 ;
        RECT 705.675 2.555 706.005 2.885 ;
        RECT 705.675 1.195 706.005 1.525 ;
        RECT 705.675 -0.165 706.005 0.165 ;
        RECT 705.68 -8.32 706 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 707.035 10.715 707.365 11.045 ;
        RECT 707.035 9.355 707.365 9.685 ;
        RECT 707.035 7.995 707.365 8.325 ;
        RECT 707.035 6.635 707.365 6.965 ;
        RECT 707.035 5.275 707.365 5.605 ;
        RECT 707.035 3.915 707.365 4.245 ;
        RECT 707.035 2.555 707.365 2.885 ;
        RECT 707.035 1.195 707.365 1.525 ;
        RECT 707.035 -0.165 707.365 0.165 ;
        RECT 707.04 -8.32 707.36 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 708.395 10.715 708.725 11.045 ;
        RECT 708.395 9.355 708.725 9.685 ;
        RECT 708.395 7.995 708.725 8.325 ;
        RECT 708.395 6.635 708.725 6.965 ;
        RECT 708.395 5.275 708.725 5.605 ;
        RECT 708.395 3.915 708.725 4.245 ;
        RECT 708.395 2.555 708.725 2.885 ;
        RECT 708.395 1.195 708.725 1.525 ;
        RECT 708.395 -0.165 708.725 0.165 ;
        RECT 708.4 -8.32 708.72 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 709.755 10.715 710.085 11.045 ;
        RECT 709.755 9.355 710.085 9.685 ;
        RECT 709.755 7.995 710.085 8.325 ;
        RECT 709.755 6.635 710.085 6.965 ;
        RECT 709.755 5.275 710.085 5.605 ;
        RECT 709.755 3.915 710.085 4.245 ;
        RECT 709.755 2.555 710.085 2.885 ;
        RECT 709.755 1.195 710.085 1.525 ;
        RECT 709.755 -0.165 710.085 0.165 ;
        RECT 709.76 -8.32 710.08 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 711.115 10.715 711.445 11.045 ;
        RECT 711.115 9.355 711.445 9.685 ;
        RECT 711.115 7.995 711.445 8.325 ;
        RECT 711.115 6.635 711.445 6.965 ;
        RECT 711.115 5.275 711.445 5.605 ;
        RECT 711.115 3.915 711.445 4.245 ;
        RECT 711.115 2.555 711.445 2.885 ;
        RECT 711.115 1.195 711.445 1.525 ;
        RECT 711.115 -0.165 711.445 0.165 ;
        RECT 711.12 -8.32 711.44 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 712.475 10.715 712.805 11.045 ;
        RECT 712.475 9.355 712.805 9.685 ;
        RECT 712.475 7.995 712.805 8.325 ;
        RECT 712.475 6.635 712.805 6.965 ;
        RECT 712.475 5.275 712.805 5.605 ;
        RECT 712.475 3.915 712.805 4.245 ;
        RECT 712.475 2.555 712.805 2.885 ;
        RECT 712.475 1.195 712.805 1.525 ;
        RECT 712.475 -0.165 712.805 0.165 ;
        RECT 712.48 -8.32 712.8 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 713.835 10.715 714.165 11.045 ;
        RECT 713.835 9.355 714.165 9.685 ;
        RECT 713.835 7.995 714.165 8.325 ;
        RECT 713.835 6.635 714.165 6.965 ;
        RECT 713.835 5.275 714.165 5.605 ;
        RECT 713.835 3.915 714.165 4.245 ;
        RECT 713.835 2.555 714.165 2.885 ;
        RECT 713.835 1.195 714.165 1.525 ;
        RECT 713.835 -0.165 714.165 0.165 ;
        RECT 713.84 -8.32 714.16 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 715.195 10.715 715.525 11.045 ;
        RECT 715.195 9.355 715.525 9.685 ;
        RECT 715.195 7.995 715.525 8.325 ;
        RECT 715.195 6.635 715.525 6.965 ;
        RECT 715.195 5.275 715.525 5.605 ;
        RECT 715.195 3.915 715.525 4.245 ;
        RECT 715.195 2.555 715.525 2.885 ;
        RECT 715.195 1.195 715.525 1.525 ;
        RECT 715.195 -0.165 715.525 0.165 ;
        RECT 715.2 -8.32 715.52 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 716.555 10.715 716.885 11.045 ;
        RECT 716.555 9.355 716.885 9.685 ;
        RECT 716.555 7.995 716.885 8.325 ;
        RECT 716.555 6.635 716.885 6.965 ;
        RECT 716.555 5.275 716.885 5.605 ;
        RECT 716.555 3.915 716.885 4.245 ;
        RECT 716.555 2.555 716.885 2.885 ;
        RECT 716.555 1.195 716.885 1.525 ;
        RECT 716.555 -0.165 716.885 0.165 ;
        RECT 716.56 -8.32 716.88 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 717.915 10.715 718.245 11.045 ;
        RECT 717.915 9.355 718.245 9.685 ;
        RECT 717.915 7.995 718.245 8.325 ;
        RECT 717.915 6.635 718.245 6.965 ;
        RECT 717.915 5.275 718.245 5.605 ;
        RECT 717.915 3.915 718.245 4.245 ;
        RECT 717.915 2.555 718.245 2.885 ;
        RECT 717.915 1.195 718.245 1.525 ;
        RECT 717.915 -0.165 718.245 0.165 ;
        RECT 717.92 -8.32 718.24 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 719.275 10.715 719.605 11.045 ;
        RECT 719.275 9.355 719.605 9.685 ;
        RECT 719.275 7.995 719.605 8.325 ;
        RECT 719.275 6.635 719.605 6.965 ;
        RECT 719.275 5.275 719.605 5.605 ;
        RECT 719.275 3.915 719.605 4.245 ;
        RECT 719.275 2.555 719.605 2.885 ;
        RECT 719.275 1.195 719.605 1.525 ;
        RECT 719.275 -0.165 719.605 0.165 ;
        RECT 719.28 -8.32 719.6 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 720.635 10.715 720.965 11.045 ;
        RECT 720.635 9.355 720.965 9.685 ;
        RECT 720.635 7.995 720.965 8.325 ;
        RECT 720.635 6.635 720.965 6.965 ;
        RECT 720.635 5.275 720.965 5.605 ;
        RECT 720.635 3.915 720.965 4.245 ;
        RECT 720.635 2.555 720.965 2.885 ;
        RECT 720.635 1.195 720.965 1.525 ;
        RECT 720.635 -0.165 720.965 0.165 ;
        RECT 720.64 -8.32 720.96 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 721.995 10.715 722.325 11.045 ;
        RECT 721.995 9.355 722.325 9.685 ;
        RECT 721.995 7.995 722.325 8.325 ;
        RECT 721.995 6.635 722.325 6.965 ;
        RECT 721.995 5.275 722.325 5.605 ;
        RECT 721.995 3.915 722.325 4.245 ;
        RECT 721.995 2.555 722.325 2.885 ;
        RECT 721.995 1.195 722.325 1.525 ;
        RECT 721.995 -0.165 722.325 0.165 ;
        RECT 722 -8.32 722.32 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 723.355 10.715 723.685 11.045 ;
        RECT 723.355 9.355 723.685 9.685 ;
        RECT 723.355 7.995 723.685 8.325 ;
        RECT 723.355 6.635 723.685 6.965 ;
        RECT 723.355 5.275 723.685 5.605 ;
        RECT 723.355 3.915 723.685 4.245 ;
        RECT 723.355 2.555 723.685 2.885 ;
        RECT 723.355 1.195 723.685 1.525 ;
        RECT 723.355 -0.165 723.685 0.165 ;
        RECT 723.36 -8.32 723.68 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 724.715 10.715 725.045 11.045 ;
        RECT 724.715 9.355 725.045 9.685 ;
        RECT 724.715 7.995 725.045 8.325 ;
        RECT 724.715 6.635 725.045 6.965 ;
        RECT 724.715 5.275 725.045 5.605 ;
        RECT 724.715 3.915 725.045 4.245 ;
        RECT 724.715 2.555 725.045 2.885 ;
        RECT 724.715 1.195 725.045 1.525 ;
        RECT 724.715 -0.165 725.045 0.165 ;
        RECT 724.72 -8.32 725.04 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 726.075 10.715 726.405 11.045 ;
        RECT 726.075 9.355 726.405 9.685 ;
        RECT 726.075 7.995 726.405 8.325 ;
        RECT 726.075 6.635 726.405 6.965 ;
        RECT 726.075 5.275 726.405 5.605 ;
        RECT 726.075 3.915 726.405 4.245 ;
        RECT 726.075 2.555 726.405 2.885 ;
        RECT 726.075 1.195 726.405 1.525 ;
        RECT 726.075 -0.165 726.405 0.165 ;
        RECT 726.08 -8.32 726.4 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 727.435 10.715 727.765 11.045 ;
        RECT 727.435 9.355 727.765 9.685 ;
        RECT 727.435 7.995 727.765 8.325 ;
        RECT 727.435 6.635 727.765 6.965 ;
        RECT 727.435 5.275 727.765 5.605 ;
        RECT 727.435 3.915 727.765 4.245 ;
        RECT 727.435 2.555 727.765 2.885 ;
        RECT 727.435 1.195 727.765 1.525 ;
        RECT 727.435 -0.165 727.765 0.165 ;
        RECT 727.44 -8.32 727.76 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 728.795 10.715 729.125 11.045 ;
        RECT 728.795 9.355 729.125 9.685 ;
        RECT 728.795 7.995 729.125 8.325 ;
        RECT 728.795 6.635 729.125 6.965 ;
        RECT 728.795 5.275 729.125 5.605 ;
        RECT 728.795 3.915 729.125 4.245 ;
        RECT 728.795 2.555 729.125 2.885 ;
        RECT 728.795 1.195 729.125 1.525 ;
        RECT 728.795 -0.165 729.125 0.165 ;
        RECT 728.8 -8.32 729.12 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 730.155 10.715 730.485 11.045 ;
        RECT 730.155 9.355 730.485 9.685 ;
        RECT 730.155 7.995 730.485 8.325 ;
        RECT 730.155 6.635 730.485 6.965 ;
        RECT 730.155 5.275 730.485 5.605 ;
        RECT 730.155 3.915 730.485 4.245 ;
        RECT 730.155 2.555 730.485 2.885 ;
        RECT 730.155 1.195 730.485 1.525 ;
        RECT 730.155 -0.165 730.485 0.165 ;
        RECT 730.16 -8.32 730.48 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 731.515 10.715 731.845 11.045 ;
        RECT 731.515 9.355 731.845 9.685 ;
        RECT 731.515 7.995 731.845 8.325 ;
        RECT 731.515 6.635 731.845 6.965 ;
        RECT 731.515 5.275 731.845 5.605 ;
        RECT 731.515 3.915 731.845 4.245 ;
        RECT 731.515 2.555 731.845 2.885 ;
        RECT 731.515 1.195 731.845 1.525 ;
        RECT 731.515 -0.165 731.845 0.165 ;
        RECT 731.52 -8.32 731.84 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 732.875 10.715 733.205 11.045 ;
        RECT 732.875 9.355 733.205 9.685 ;
        RECT 732.875 7.995 733.205 8.325 ;
        RECT 732.875 6.635 733.205 6.965 ;
        RECT 732.875 5.275 733.205 5.605 ;
        RECT 732.875 3.915 733.205 4.245 ;
        RECT 732.875 2.555 733.205 2.885 ;
        RECT 732.875 1.195 733.205 1.525 ;
        RECT 732.875 -0.165 733.205 0.165 ;
        RECT 732.88 -8.32 733.2 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 734.235 10.715 734.565 11.045 ;
        RECT 734.235 9.355 734.565 9.685 ;
        RECT 734.235 7.995 734.565 8.325 ;
        RECT 734.235 6.635 734.565 6.965 ;
        RECT 734.235 5.275 734.565 5.605 ;
        RECT 734.235 3.915 734.565 4.245 ;
        RECT 734.235 2.555 734.565 2.885 ;
        RECT 734.235 1.195 734.565 1.525 ;
        RECT 734.235 -0.165 734.565 0.165 ;
        RECT 734.24 -8.32 734.56 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 735.595 10.715 735.925 11.045 ;
        RECT 735.595 9.355 735.925 9.685 ;
        RECT 735.595 7.995 735.925 8.325 ;
        RECT 735.595 6.635 735.925 6.965 ;
        RECT 735.595 5.275 735.925 5.605 ;
        RECT 735.595 3.915 735.925 4.245 ;
        RECT 735.595 2.555 735.925 2.885 ;
        RECT 735.595 1.195 735.925 1.525 ;
        RECT 735.595 -0.165 735.925 0.165 ;
        RECT 735.6 -8.32 735.92 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 736.955 10.715 737.285 11.045 ;
        RECT 736.955 9.355 737.285 9.685 ;
        RECT 736.955 7.995 737.285 8.325 ;
        RECT 736.955 6.635 737.285 6.965 ;
        RECT 736.955 5.275 737.285 5.605 ;
        RECT 736.955 3.915 737.285 4.245 ;
        RECT 736.955 2.555 737.285 2.885 ;
        RECT 736.955 1.195 737.285 1.525 ;
        RECT 736.955 -0.165 737.285 0.165 ;
        RECT 736.96 -8.32 737.28 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 738.315 10.715 738.645 11.045 ;
        RECT 738.315 9.355 738.645 9.685 ;
        RECT 738.315 7.995 738.645 8.325 ;
        RECT 738.315 6.635 738.645 6.965 ;
        RECT 738.315 5.275 738.645 5.605 ;
        RECT 738.315 3.915 738.645 4.245 ;
        RECT 738.315 2.555 738.645 2.885 ;
        RECT 738.315 1.195 738.645 1.525 ;
        RECT 738.315 -0.165 738.645 0.165 ;
        RECT 738.32 -8.32 738.64 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 739.675 10.715 740.005 11.045 ;
        RECT 739.675 9.355 740.005 9.685 ;
        RECT 739.675 7.995 740.005 8.325 ;
        RECT 739.675 6.635 740.005 6.965 ;
        RECT 739.675 5.275 740.005 5.605 ;
        RECT 739.675 3.915 740.005 4.245 ;
        RECT 739.675 2.555 740.005 2.885 ;
        RECT 739.675 1.195 740.005 1.525 ;
        RECT 739.675 -0.165 740.005 0.165 ;
        RECT 739.68 -8.32 740 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 741.035 10.715 741.365 11.045 ;
        RECT 741.035 9.355 741.365 9.685 ;
        RECT 741.035 7.995 741.365 8.325 ;
        RECT 741.035 6.635 741.365 6.965 ;
        RECT 741.035 5.275 741.365 5.605 ;
        RECT 741.035 3.915 741.365 4.245 ;
        RECT 741.035 2.555 741.365 2.885 ;
        RECT 741.035 1.195 741.365 1.525 ;
        RECT 741.035 -0.165 741.365 0.165 ;
        RECT 741.04 -8.32 741.36 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 742.395 10.715 742.725 11.045 ;
        RECT 742.395 9.355 742.725 9.685 ;
        RECT 742.395 7.995 742.725 8.325 ;
        RECT 742.395 6.635 742.725 6.965 ;
        RECT 742.395 5.275 742.725 5.605 ;
        RECT 742.395 3.915 742.725 4.245 ;
        RECT 742.395 2.555 742.725 2.885 ;
        RECT 742.395 1.195 742.725 1.525 ;
        RECT 742.395 -0.165 742.725 0.165 ;
        RECT 742.4 -8.32 742.72 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 743.755 10.715 744.085 11.045 ;
        RECT 743.755 9.355 744.085 9.685 ;
        RECT 743.755 7.995 744.085 8.325 ;
        RECT 743.755 6.635 744.085 6.965 ;
        RECT 743.755 5.275 744.085 5.605 ;
        RECT 743.755 3.915 744.085 4.245 ;
        RECT 743.755 2.555 744.085 2.885 ;
        RECT 743.755 1.195 744.085 1.525 ;
        RECT 743.755 -0.165 744.085 0.165 ;
        RECT 743.76 -8.32 744.08 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 745.115 10.715 745.445 11.045 ;
        RECT 745.115 9.355 745.445 9.685 ;
        RECT 745.115 7.995 745.445 8.325 ;
        RECT 745.115 6.635 745.445 6.965 ;
        RECT 745.115 5.275 745.445 5.605 ;
        RECT 745.115 3.915 745.445 4.245 ;
        RECT 745.115 2.555 745.445 2.885 ;
        RECT 745.115 1.195 745.445 1.525 ;
        RECT 745.115 -0.165 745.445 0.165 ;
        RECT 745.12 -8.32 745.44 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 746.475 10.715 746.805 11.045 ;
        RECT 746.475 9.355 746.805 9.685 ;
        RECT 746.475 7.995 746.805 8.325 ;
        RECT 746.475 6.635 746.805 6.965 ;
        RECT 746.475 5.275 746.805 5.605 ;
        RECT 746.475 3.915 746.805 4.245 ;
        RECT 746.475 2.555 746.805 2.885 ;
        RECT 746.475 1.195 746.805 1.525 ;
        RECT 746.475 -0.165 746.805 0.165 ;
        RECT 746.48 -8.32 746.8 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 747.835 10.715 748.165 11.045 ;
        RECT 747.835 9.355 748.165 9.685 ;
        RECT 747.835 7.995 748.165 8.325 ;
        RECT 747.835 6.635 748.165 6.965 ;
        RECT 747.835 5.275 748.165 5.605 ;
        RECT 747.835 3.915 748.165 4.245 ;
        RECT 747.835 2.555 748.165 2.885 ;
        RECT 747.835 1.195 748.165 1.525 ;
        RECT 747.835 -0.165 748.165 0.165 ;
        RECT 747.84 -8.32 748.16 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 749.195 10.715 749.525 11.045 ;
        RECT 749.195 9.355 749.525 9.685 ;
        RECT 749.195 7.995 749.525 8.325 ;
        RECT 749.195 6.635 749.525 6.965 ;
        RECT 749.195 5.275 749.525 5.605 ;
        RECT 749.195 3.915 749.525 4.245 ;
        RECT 749.195 2.555 749.525 2.885 ;
        RECT 749.195 1.195 749.525 1.525 ;
        RECT 749.195 -0.165 749.525 0.165 ;
        RECT 749.2 -8.32 749.52 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 750.555 10.715 750.885 11.045 ;
        RECT 750.555 9.355 750.885 9.685 ;
        RECT 750.555 7.995 750.885 8.325 ;
        RECT 750.555 6.635 750.885 6.965 ;
        RECT 750.555 5.275 750.885 5.605 ;
        RECT 750.555 3.915 750.885 4.245 ;
        RECT 750.555 2.555 750.885 2.885 ;
        RECT 750.555 1.195 750.885 1.525 ;
        RECT 750.555 -0.165 750.885 0.165 ;
        RECT 750.56 -8.32 750.88 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 751.915 10.715 752.245 11.045 ;
        RECT 751.915 9.355 752.245 9.685 ;
        RECT 751.915 7.995 752.245 8.325 ;
        RECT 751.915 6.635 752.245 6.965 ;
        RECT 751.915 5.275 752.245 5.605 ;
        RECT 751.915 3.915 752.245 4.245 ;
        RECT 751.915 2.555 752.245 2.885 ;
        RECT 751.915 1.195 752.245 1.525 ;
        RECT 751.915 -0.165 752.245 0.165 ;
        RECT 751.92 -8.32 752.24 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 753.275 10.715 753.605 11.045 ;
        RECT 753.275 9.355 753.605 9.685 ;
        RECT 753.275 7.995 753.605 8.325 ;
        RECT 753.275 6.635 753.605 6.965 ;
        RECT 753.275 5.275 753.605 5.605 ;
        RECT 753.275 3.915 753.605 4.245 ;
        RECT 753.275 2.555 753.605 2.885 ;
        RECT 753.275 1.195 753.605 1.525 ;
        RECT 753.275 -0.165 753.605 0.165 ;
        RECT 753.28 -8.32 753.6 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 754.635 10.715 754.965 11.045 ;
        RECT 754.635 9.355 754.965 9.685 ;
        RECT 754.635 7.995 754.965 8.325 ;
        RECT 754.635 6.635 754.965 6.965 ;
        RECT 754.635 5.275 754.965 5.605 ;
        RECT 754.635 3.915 754.965 4.245 ;
        RECT 754.635 2.555 754.965 2.885 ;
        RECT 754.635 1.195 754.965 1.525 ;
        RECT 754.635 -0.165 754.965 0.165 ;
        RECT 754.64 -8.32 754.96 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 755.995 10.715 756.325 11.045 ;
        RECT 755.995 9.355 756.325 9.685 ;
        RECT 755.995 7.995 756.325 8.325 ;
        RECT 755.995 6.635 756.325 6.965 ;
        RECT 755.995 5.275 756.325 5.605 ;
        RECT 755.995 3.915 756.325 4.245 ;
        RECT 755.995 2.555 756.325 2.885 ;
        RECT 755.995 1.195 756.325 1.525 ;
        RECT 755.995 -0.165 756.325 0.165 ;
        RECT 756 -8.32 756.32 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 757.355 10.715 757.685 11.045 ;
        RECT 757.355 9.355 757.685 9.685 ;
        RECT 757.355 7.995 757.685 8.325 ;
        RECT 757.355 6.635 757.685 6.965 ;
        RECT 757.355 5.275 757.685 5.605 ;
        RECT 757.355 3.915 757.685 4.245 ;
        RECT 757.355 2.555 757.685 2.885 ;
        RECT 757.355 1.195 757.685 1.525 ;
        RECT 757.355 -0.165 757.685 0.165 ;
        RECT 757.36 -8.32 757.68 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 758.715 10.715 759.045 11.045 ;
        RECT 758.715 9.355 759.045 9.685 ;
        RECT 758.715 7.995 759.045 8.325 ;
        RECT 758.715 6.635 759.045 6.965 ;
        RECT 758.715 5.275 759.045 5.605 ;
        RECT 758.715 3.915 759.045 4.245 ;
        RECT 758.715 2.555 759.045 2.885 ;
        RECT 758.715 1.195 759.045 1.525 ;
        RECT 758.715 -0.165 759.045 0.165 ;
        RECT 758.72 -8.32 759.04 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 760.075 10.715 760.405 11.045 ;
        RECT 760.075 9.355 760.405 9.685 ;
        RECT 760.075 7.995 760.405 8.325 ;
        RECT 760.075 6.635 760.405 6.965 ;
        RECT 760.075 5.275 760.405 5.605 ;
        RECT 760.075 3.915 760.405 4.245 ;
        RECT 760.075 2.555 760.405 2.885 ;
        RECT 760.075 1.195 760.405 1.525 ;
        RECT 760.075 -0.165 760.405 0.165 ;
        RECT 760.08 -8.32 760.4 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 761.435 10.715 761.765 11.045 ;
        RECT 761.435 9.355 761.765 9.685 ;
        RECT 761.435 7.995 761.765 8.325 ;
        RECT 761.435 6.635 761.765 6.965 ;
        RECT 761.435 5.275 761.765 5.605 ;
        RECT 761.435 3.915 761.765 4.245 ;
        RECT 761.435 2.555 761.765 2.885 ;
        RECT 761.435 1.195 761.765 1.525 ;
        RECT 761.435 -0.165 761.765 0.165 ;
        RECT 761.44 -8.32 761.76 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 762.795 13.435 763.125 13.765 ;
        RECT 762.795 10.715 763.125 11.045 ;
        RECT 762.795 9.355 763.125 9.685 ;
        RECT 762.795 7.995 763.125 8.325 ;
        RECT 762.795 6.635 763.125 6.965 ;
        RECT 762.795 5.275 763.125 5.605 ;
        RECT 762.795 3.915 763.125 4.245 ;
        RECT 762.795 2.555 763.125 2.885 ;
        RECT 762.795 1.195 763.125 1.525 ;
        RECT 762.795 -0.165 763.125 0.165 ;
        RECT 762.8 -8.32 763.12 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 764.155 13.435 764.485 13.765 ;
        RECT 764.155 10.715 764.485 11.045 ;
        RECT 764.155 9.355 764.485 9.685 ;
        RECT 764.155 7.995 764.485 8.325 ;
        RECT 764.155 6.635 764.485 6.965 ;
        RECT 764.155 5.275 764.485 5.605 ;
        RECT 764.155 3.915 764.485 4.245 ;
        RECT 764.155 2.555 764.485 2.885 ;
        RECT 764.155 1.195 764.485 1.525 ;
        RECT 764.155 -0.165 764.485 0.165 ;
        RECT 764.16 -8.32 764.48 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 765.515 13.435 765.845 13.765 ;
        RECT 765.515 12.075 765.845 12.405 ;
        RECT 765.515 10.715 765.845 11.045 ;
        RECT 765.515 9.355 765.845 9.685 ;
        RECT 765.515 7.995 765.845 8.325 ;
        RECT 765.515 6.635 765.845 6.965 ;
        RECT 765.515 5.275 765.845 5.605 ;
        RECT 765.515 3.915 765.845 4.245 ;
        RECT 765.515 2.555 765.845 2.885 ;
        RECT 765.515 1.195 765.845 1.525 ;
        RECT 765.515 -0.165 765.845 0.165 ;
        RECT 765.52 -8.32 765.84 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 766.875 13.435 767.205 13.765 ;
        RECT 766.875 12.075 767.205 12.405 ;
        RECT 766.875 10.715 767.205 11.045 ;
        RECT 766.875 9.355 767.205 9.685 ;
        RECT 766.875 7.995 767.205 8.325 ;
        RECT 766.875 6.635 767.205 6.965 ;
        RECT 766.875 5.275 767.205 5.605 ;
        RECT 766.875 3.915 767.205 4.245 ;
        RECT 766.875 2.555 767.205 2.885 ;
        RECT 766.875 1.195 767.205 1.525 ;
        RECT 766.875 -0.165 767.205 0.165 ;
        RECT 766.88 -8.32 767.2 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 768.235 14.795 768.565 15.125 ;
        RECT 768.235 13.435 768.565 13.765 ;
        RECT 768.235 12.075 768.565 12.405 ;
        RECT 768.235 10.715 768.565 11.045 ;
        RECT 768.235 9.355 768.565 9.685 ;
        RECT 768.235 7.995 768.565 8.325 ;
        RECT 768.235 6.635 768.565 6.965 ;
        RECT 768.235 5.275 768.565 5.605 ;
        RECT 768.235 3.915 768.565 4.245 ;
        RECT 768.235 2.555 768.565 2.885 ;
        RECT 768.235 1.195 768.565 1.525 ;
        RECT 768.235 -0.165 768.565 0.165 ;
        RECT 768.24 -8.32 768.56 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 498.955 10.715 499.285 11.045 ;
        RECT 498.955 9.355 499.285 9.685 ;
        RECT 498.955 7.995 499.285 8.325 ;
        RECT 498.955 6.635 499.285 6.965 ;
        RECT 498.955 5.275 499.285 5.605 ;
        RECT 498.955 3.915 499.285 4.245 ;
        RECT 498.955 2.555 499.285 2.885 ;
        RECT 498.955 1.195 499.285 1.525 ;
        RECT 498.955 -0.165 499.285 0.165 ;
        RECT 498.96 -8.32 499.28 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 500.315 10.715 500.645 11.045 ;
        RECT 500.315 9.355 500.645 9.685 ;
        RECT 500.315 7.995 500.645 8.325 ;
        RECT 500.315 6.635 500.645 6.965 ;
        RECT 500.315 5.275 500.645 5.605 ;
        RECT 500.315 3.915 500.645 4.245 ;
        RECT 500.315 2.555 500.645 2.885 ;
        RECT 500.315 1.195 500.645 1.525 ;
        RECT 500.315 -0.165 500.645 0.165 ;
        RECT 500.32 -8.32 500.64 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 501.675 10.715 502.005 11.045 ;
        RECT 501.675 9.355 502.005 9.685 ;
        RECT 501.675 7.995 502.005 8.325 ;
        RECT 501.675 6.635 502.005 6.965 ;
        RECT 501.675 5.275 502.005 5.605 ;
        RECT 501.675 3.915 502.005 4.245 ;
        RECT 501.675 2.555 502.005 2.885 ;
        RECT 501.675 1.195 502.005 1.525 ;
        RECT 501.675 -0.165 502.005 0.165 ;
        RECT 501.68 -8.32 502 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 503.035 10.715 503.365 11.045 ;
        RECT 503.035 9.355 503.365 9.685 ;
        RECT 503.035 7.995 503.365 8.325 ;
        RECT 503.035 6.635 503.365 6.965 ;
        RECT 503.035 5.275 503.365 5.605 ;
        RECT 503.035 3.915 503.365 4.245 ;
        RECT 503.035 2.555 503.365 2.885 ;
        RECT 503.035 1.195 503.365 1.525 ;
        RECT 503.035 -0.165 503.365 0.165 ;
        RECT 503.04 -8.32 503.36 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 504.395 10.715 504.725 11.045 ;
        RECT 504.395 9.355 504.725 9.685 ;
        RECT 504.395 7.995 504.725 8.325 ;
        RECT 504.395 6.635 504.725 6.965 ;
        RECT 504.395 5.275 504.725 5.605 ;
        RECT 504.395 3.915 504.725 4.245 ;
        RECT 504.395 2.555 504.725 2.885 ;
        RECT 504.395 1.195 504.725 1.525 ;
        RECT 504.395 -0.165 504.725 0.165 ;
        RECT 504.4 -8.32 504.72 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 505.755 10.715 506.085 11.045 ;
        RECT 505.755 9.355 506.085 9.685 ;
        RECT 505.755 7.995 506.085 8.325 ;
        RECT 505.755 6.635 506.085 6.965 ;
        RECT 505.755 5.275 506.085 5.605 ;
        RECT 505.755 3.915 506.085 4.245 ;
        RECT 505.755 2.555 506.085 2.885 ;
        RECT 505.755 1.195 506.085 1.525 ;
        RECT 505.755 -0.165 506.085 0.165 ;
        RECT 505.76 -8.32 506.08 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 507.115 10.715 507.445 11.045 ;
        RECT 507.115 9.355 507.445 9.685 ;
        RECT 507.115 7.995 507.445 8.325 ;
        RECT 507.115 6.635 507.445 6.965 ;
        RECT 507.115 5.275 507.445 5.605 ;
        RECT 507.115 3.915 507.445 4.245 ;
        RECT 507.115 2.555 507.445 2.885 ;
        RECT 507.115 1.195 507.445 1.525 ;
        RECT 507.115 -0.165 507.445 0.165 ;
        RECT 507.12 -8.32 507.44 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 508.475 10.715 508.805 11.045 ;
        RECT 508.475 9.355 508.805 9.685 ;
        RECT 508.475 7.995 508.805 8.325 ;
        RECT 508.475 6.635 508.805 6.965 ;
        RECT 508.475 5.275 508.805 5.605 ;
        RECT 508.475 3.915 508.805 4.245 ;
        RECT 508.475 2.555 508.805 2.885 ;
        RECT 508.475 1.195 508.805 1.525 ;
        RECT 508.475 -0.165 508.805 0.165 ;
        RECT 508.48 -8.32 508.8 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 509.835 10.715 510.165 11.045 ;
        RECT 509.835 9.355 510.165 9.685 ;
        RECT 509.835 7.995 510.165 8.325 ;
        RECT 509.835 6.635 510.165 6.965 ;
        RECT 509.835 5.275 510.165 5.605 ;
        RECT 509.835 3.915 510.165 4.245 ;
        RECT 509.835 2.555 510.165 2.885 ;
        RECT 509.835 1.195 510.165 1.525 ;
        RECT 509.835 -0.165 510.165 0.165 ;
        RECT 509.84 -8.32 510.16 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 511.195 10.715 511.525 11.045 ;
        RECT 511.195 9.355 511.525 9.685 ;
        RECT 511.195 7.995 511.525 8.325 ;
        RECT 511.195 6.635 511.525 6.965 ;
        RECT 511.195 5.275 511.525 5.605 ;
        RECT 511.195 3.915 511.525 4.245 ;
        RECT 511.195 2.555 511.525 2.885 ;
        RECT 511.195 1.195 511.525 1.525 ;
        RECT 511.195 -0.165 511.525 0.165 ;
        RECT 511.2 -8.32 511.52 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 512.555 10.715 512.885 11.045 ;
        RECT 512.555 9.355 512.885 9.685 ;
        RECT 512.555 7.995 512.885 8.325 ;
        RECT 512.555 6.635 512.885 6.965 ;
        RECT 512.555 5.275 512.885 5.605 ;
        RECT 512.555 3.915 512.885 4.245 ;
        RECT 512.555 2.555 512.885 2.885 ;
        RECT 512.555 1.195 512.885 1.525 ;
        RECT 512.555 -0.165 512.885 0.165 ;
        RECT 512.56 -8.32 512.88 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 513.915 10.715 514.245 11.045 ;
        RECT 513.915 9.355 514.245 9.685 ;
        RECT 513.915 7.995 514.245 8.325 ;
        RECT 513.915 6.635 514.245 6.965 ;
        RECT 513.915 5.275 514.245 5.605 ;
        RECT 513.915 3.915 514.245 4.245 ;
        RECT 513.915 2.555 514.245 2.885 ;
        RECT 513.915 1.195 514.245 1.525 ;
        RECT 513.915 -0.165 514.245 0.165 ;
        RECT 513.92 -8.32 514.24 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 515.275 10.715 515.605 11.045 ;
        RECT 515.275 9.355 515.605 9.685 ;
        RECT 515.275 7.995 515.605 8.325 ;
        RECT 515.275 6.635 515.605 6.965 ;
        RECT 515.275 5.275 515.605 5.605 ;
        RECT 515.275 3.915 515.605 4.245 ;
        RECT 515.275 2.555 515.605 2.885 ;
        RECT 515.275 1.195 515.605 1.525 ;
        RECT 515.275 -0.165 515.605 0.165 ;
        RECT 515.28 -8.32 515.6 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 516.635 10.715 516.965 11.045 ;
        RECT 516.635 9.355 516.965 9.685 ;
        RECT 516.635 7.995 516.965 8.325 ;
        RECT 516.635 6.635 516.965 6.965 ;
        RECT 516.635 5.275 516.965 5.605 ;
        RECT 516.635 3.915 516.965 4.245 ;
        RECT 516.635 2.555 516.965 2.885 ;
        RECT 516.635 1.195 516.965 1.525 ;
        RECT 516.635 -0.165 516.965 0.165 ;
        RECT 516.64 -8.32 516.96 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 517.995 10.715 518.325 11.045 ;
        RECT 517.995 9.355 518.325 9.685 ;
        RECT 517.995 7.995 518.325 8.325 ;
        RECT 517.995 6.635 518.325 6.965 ;
        RECT 517.995 5.275 518.325 5.605 ;
        RECT 517.995 3.915 518.325 4.245 ;
        RECT 517.995 2.555 518.325 2.885 ;
        RECT 517.995 1.195 518.325 1.525 ;
        RECT 517.995 -0.165 518.325 0.165 ;
        RECT 518 -8.32 518.32 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 519.355 10.715 519.685 11.045 ;
        RECT 519.355 9.355 519.685 9.685 ;
        RECT 519.355 7.995 519.685 8.325 ;
        RECT 519.355 6.635 519.685 6.965 ;
        RECT 519.355 5.275 519.685 5.605 ;
        RECT 519.355 3.915 519.685 4.245 ;
        RECT 519.355 2.555 519.685 2.885 ;
        RECT 519.355 1.195 519.685 1.525 ;
        RECT 519.355 -0.165 519.685 0.165 ;
        RECT 519.36 -8.32 519.68 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 520.715 10.715 521.045 11.045 ;
        RECT 520.715 9.355 521.045 9.685 ;
        RECT 520.715 7.995 521.045 8.325 ;
        RECT 520.715 6.635 521.045 6.965 ;
        RECT 520.715 5.275 521.045 5.605 ;
        RECT 520.715 3.915 521.045 4.245 ;
        RECT 520.715 2.555 521.045 2.885 ;
        RECT 520.715 1.195 521.045 1.525 ;
        RECT 520.715 -0.165 521.045 0.165 ;
        RECT 520.72 -8.32 521.04 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 522.075 10.715 522.405 11.045 ;
        RECT 522.075 9.355 522.405 9.685 ;
        RECT 522.075 7.995 522.405 8.325 ;
        RECT 522.075 6.635 522.405 6.965 ;
        RECT 522.075 5.275 522.405 5.605 ;
        RECT 522.075 3.915 522.405 4.245 ;
        RECT 522.075 2.555 522.405 2.885 ;
        RECT 522.075 1.195 522.405 1.525 ;
        RECT 522.075 -0.165 522.405 0.165 ;
        RECT 522.08 -8.32 522.4 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 523.435 10.715 523.765 11.045 ;
        RECT 523.435 9.355 523.765 9.685 ;
        RECT 523.435 7.995 523.765 8.325 ;
        RECT 523.435 6.635 523.765 6.965 ;
        RECT 523.435 5.275 523.765 5.605 ;
        RECT 523.435 3.915 523.765 4.245 ;
        RECT 523.435 2.555 523.765 2.885 ;
        RECT 523.435 1.195 523.765 1.525 ;
        RECT 523.435 -0.165 523.765 0.165 ;
        RECT 523.44 -8.32 523.76 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 524.795 10.715 525.125 11.045 ;
        RECT 524.795 9.355 525.125 9.685 ;
        RECT 524.795 7.995 525.125 8.325 ;
        RECT 524.795 6.635 525.125 6.965 ;
        RECT 524.795 5.275 525.125 5.605 ;
        RECT 524.795 3.915 525.125 4.245 ;
        RECT 524.795 2.555 525.125 2.885 ;
        RECT 524.795 1.195 525.125 1.525 ;
        RECT 524.795 -0.165 525.125 0.165 ;
        RECT 524.8 -8.32 525.12 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 526.155 10.715 526.485 11.045 ;
        RECT 526.155 9.355 526.485 9.685 ;
        RECT 526.155 7.995 526.485 8.325 ;
        RECT 526.155 6.635 526.485 6.965 ;
        RECT 526.155 5.275 526.485 5.605 ;
        RECT 526.155 3.915 526.485 4.245 ;
        RECT 526.155 2.555 526.485 2.885 ;
        RECT 526.155 1.195 526.485 1.525 ;
        RECT 526.155 -0.165 526.485 0.165 ;
        RECT 526.16 -8.32 526.48 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 527.515 10.715 527.845 11.045 ;
        RECT 527.515 9.355 527.845 9.685 ;
        RECT 527.515 7.995 527.845 8.325 ;
        RECT 527.515 6.635 527.845 6.965 ;
        RECT 527.515 5.275 527.845 5.605 ;
        RECT 527.515 3.915 527.845 4.245 ;
        RECT 527.515 2.555 527.845 2.885 ;
        RECT 527.515 1.195 527.845 1.525 ;
        RECT 527.515 -0.165 527.845 0.165 ;
        RECT 527.52 -8.32 527.84 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 528.875 10.715 529.205 11.045 ;
        RECT 528.875 9.355 529.205 9.685 ;
        RECT 528.875 7.995 529.205 8.325 ;
        RECT 528.875 6.635 529.205 6.965 ;
        RECT 528.875 5.275 529.205 5.605 ;
        RECT 528.875 3.915 529.205 4.245 ;
        RECT 528.875 2.555 529.205 2.885 ;
        RECT 528.875 1.195 529.205 1.525 ;
        RECT 528.875 -0.165 529.205 0.165 ;
        RECT 528.88 -8.32 529.2 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 530.235 10.715 530.565 11.045 ;
        RECT 530.235 9.355 530.565 9.685 ;
        RECT 530.235 7.995 530.565 8.325 ;
        RECT 530.235 6.635 530.565 6.965 ;
        RECT 530.235 5.275 530.565 5.605 ;
        RECT 530.235 3.915 530.565 4.245 ;
        RECT 530.235 2.555 530.565 2.885 ;
        RECT 530.235 1.195 530.565 1.525 ;
        RECT 530.235 -0.165 530.565 0.165 ;
        RECT 530.24 -8.32 530.56 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 531.595 10.715 531.925 11.045 ;
        RECT 531.595 9.355 531.925 9.685 ;
        RECT 531.595 7.995 531.925 8.325 ;
        RECT 531.595 6.635 531.925 6.965 ;
        RECT 531.595 5.275 531.925 5.605 ;
        RECT 531.595 3.915 531.925 4.245 ;
        RECT 531.595 2.555 531.925 2.885 ;
        RECT 531.595 1.195 531.925 1.525 ;
        RECT 531.595 -0.165 531.925 0.165 ;
        RECT 531.6 -8.32 531.92 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 532.955 10.715 533.285 11.045 ;
        RECT 532.955 9.355 533.285 9.685 ;
        RECT 532.955 7.995 533.285 8.325 ;
        RECT 532.955 6.635 533.285 6.965 ;
        RECT 532.955 5.275 533.285 5.605 ;
        RECT 532.955 3.915 533.285 4.245 ;
        RECT 532.955 2.555 533.285 2.885 ;
        RECT 532.955 1.195 533.285 1.525 ;
        RECT 532.955 -0.165 533.285 0.165 ;
        RECT 532.96 -8.32 533.28 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 534.315 10.715 534.645 11.045 ;
        RECT 534.315 9.355 534.645 9.685 ;
        RECT 534.315 7.995 534.645 8.325 ;
        RECT 534.315 6.635 534.645 6.965 ;
        RECT 534.315 5.275 534.645 5.605 ;
        RECT 534.315 3.915 534.645 4.245 ;
        RECT 534.315 2.555 534.645 2.885 ;
        RECT 534.315 1.195 534.645 1.525 ;
        RECT 534.315 -0.165 534.645 0.165 ;
        RECT 534.32 -8.32 534.64 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 535.675 10.715 536.005 11.045 ;
        RECT 535.675 9.355 536.005 9.685 ;
        RECT 535.675 7.995 536.005 8.325 ;
        RECT 535.675 6.635 536.005 6.965 ;
        RECT 535.675 5.275 536.005 5.605 ;
        RECT 535.675 3.915 536.005 4.245 ;
        RECT 535.675 2.555 536.005 2.885 ;
        RECT 535.675 1.195 536.005 1.525 ;
        RECT 535.675 -0.165 536.005 0.165 ;
        RECT 535.68 -8.32 536 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 537.035 10.715 537.365 11.045 ;
        RECT 537.035 9.355 537.365 9.685 ;
        RECT 537.035 7.995 537.365 8.325 ;
        RECT 537.035 6.635 537.365 6.965 ;
        RECT 537.035 5.275 537.365 5.605 ;
        RECT 537.035 3.915 537.365 4.245 ;
        RECT 537.035 2.555 537.365 2.885 ;
        RECT 537.035 1.195 537.365 1.525 ;
        RECT 537.035 -0.165 537.365 0.165 ;
        RECT 537.04 -8.32 537.36 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 538.395 10.715 538.725 11.045 ;
        RECT 538.395 9.355 538.725 9.685 ;
        RECT 538.395 7.995 538.725 8.325 ;
        RECT 538.395 6.635 538.725 6.965 ;
        RECT 538.395 5.275 538.725 5.605 ;
        RECT 538.395 3.915 538.725 4.245 ;
        RECT 538.395 2.555 538.725 2.885 ;
        RECT 538.395 1.195 538.725 1.525 ;
        RECT 538.395 -0.165 538.725 0.165 ;
        RECT 538.4 -8.32 538.72 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 539.755 10.715 540.085 11.045 ;
        RECT 539.755 9.355 540.085 9.685 ;
        RECT 539.755 7.995 540.085 8.325 ;
        RECT 539.755 6.635 540.085 6.965 ;
        RECT 539.755 5.275 540.085 5.605 ;
        RECT 539.755 3.915 540.085 4.245 ;
        RECT 539.755 2.555 540.085 2.885 ;
        RECT 539.755 1.195 540.085 1.525 ;
        RECT 539.755 -0.165 540.085 0.165 ;
        RECT 539.76 -8.32 540.08 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 541.115 10.715 541.445 11.045 ;
        RECT 541.115 9.355 541.445 9.685 ;
        RECT 541.115 7.995 541.445 8.325 ;
        RECT 541.115 6.635 541.445 6.965 ;
        RECT 541.115 5.275 541.445 5.605 ;
        RECT 541.115 3.915 541.445 4.245 ;
        RECT 541.115 2.555 541.445 2.885 ;
        RECT 541.115 1.195 541.445 1.525 ;
        RECT 541.115 -0.165 541.445 0.165 ;
        RECT 541.12 -8.32 541.44 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 542.475 10.715 542.805 11.045 ;
        RECT 542.475 9.355 542.805 9.685 ;
        RECT 542.475 7.995 542.805 8.325 ;
        RECT 542.475 6.635 542.805 6.965 ;
        RECT 542.475 5.275 542.805 5.605 ;
        RECT 542.475 3.915 542.805 4.245 ;
        RECT 542.475 2.555 542.805 2.885 ;
        RECT 542.475 1.195 542.805 1.525 ;
        RECT 542.475 -0.165 542.805 0.165 ;
        RECT 542.48 -8.32 542.8 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 543.835 10.715 544.165 11.045 ;
        RECT 543.835 9.355 544.165 9.685 ;
        RECT 543.835 7.995 544.165 8.325 ;
        RECT 543.835 6.635 544.165 6.965 ;
        RECT 543.835 5.275 544.165 5.605 ;
        RECT 543.835 3.915 544.165 4.245 ;
        RECT 543.835 2.555 544.165 2.885 ;
        RECT 543.835 1.195 544.165 1.525 ;
        RECT 543.835 -0.165 544.165 0.165 ;
        RECT 543.84 -8.32 544.16 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 545.195 10.715 545.525 11.045 ;
        RECT 545.195 9.355 545.525 9.685 ;
        RECT 545.195 7.995 545.525 8.325 ;
        RECT 545.195 6.635 545.525 6.965 ;
        RECT 545.195 5.275 545.525 5.605 ;
        RECT 545.195 3.915 545.525 4.245 ;
        RECT 545.195 2.555 545.525 2.885 ;
        RECT 545.195 1.195 545.525 1.525 ;
        RECT 545.195 -0.165 545.525 0.165 ;
        RECT 545.2 -8.32 545.52 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 546.555 10.715 546.885 11.045 ;
        RECT 546.555 9.355 546.885 9.685 ;
        RECT 546.555 7.995 546.885 8.325 ;
        RECT 546.555 6.635 546.885 6.965 ;
        RECT 546.555 5.275 546.885 5.605 ;
        RECT 546.555 3.915 546.885 4.245 ;
        RECT 546.555 2.555 546.885 2.885 ;
        RECT 546.555 1.195 546.885 1.525 ;
        RECT 546.555 -0.165 546.885 0.165 ;
        RECT 546.56 -8.32 546.88 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 547.915 10.715 548.245 11.045 ;
        RECT 547.915 9.355 548.245 9.685 ;
        RECT 547.915 7.995 548.245 8.325 ;
        RECT 547.915 6.635 548.245 6.965 ;
        RECT 547.915 5.275 548.245 5.605 ;
        RECT 547.915 3.915 548.245 4.245 ;
        RECT 547.915 2.555 548.245 2.885 ;
        RECT 547.915 1.195 548.245 1.525 ;
        RECT 547.915 -0.165 548.245 0.165 ;
        RECT 547.92 -8.32 548.24 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 549.275 10.715 549.605 11.045 ;
        RECT 549.275 9.355 549.605 9.685 ;
        RECT 549.275 7.995 549.605 8.325 ;
        RECT 549.275 6.635 549.605 6.965 ;
        RECT 549.275 5.275 549.605 5.605 ;
        RECT 549.275 3.915 549.605 4.245 ;
        RECT 549.275 2.555 549.605 2.885 ;
        RECT 549.275 1.195 549.605 1.525 ;
        RECT 549.275 -0.165 549.605 0.165 ;
        RECT 549.28 -8.32 549.6 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 550.635 10.715 550.965 11.045 ;
        RECT 550.635 9.355 550.965 9.685 ;
        RECT 550.635 7.995 550.965 8.325 ;
        RECT 550.635 6.635 550.965 6.965 ;
        RECT 550.635 5.275 550.965 5.605 ;
        RECT 550.635 3.915 550.965 4.245 ;
        RECT 550.635 2.555 550.965 2.885 ;
        RECT 550.635 1.195 550.965 1.525 ;
        RECT 550.635 -0.165 550.965 0.165 ;
        RECT 550.64 -8.32 550.96 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 551.995 10.715 552.325 11.045 ;
        RECT 551.995 9.355 552.325 9.685 ;
        RECT 551.995 7.995 552.325 8.325 ;
        RECT 551.995 6.635 552.325 6.965 ;
        RECT 551.995 5.275 552.325 5.605 ;
        RECT 551.995 3.915 552.325 4.245 ;
        RECT 551.995 2.555 552.325 2.885 ;
        RECT 551.995 1.195 552.325 1.525 ;
        RECT 551.995 -0.165 552.325 0.165 ;
        RECT 552 -8.32 552.32 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 553.355 10.715 553.685 11.045 ;
        RECT 553.355 9.355 553.685 9.685 ;
        RECT 553.355 7.995 553.685 8.325 ;
        RECT 553.355 6.635 553.685 6.965 ;
        RECT 553.355 5.275 553.685 5.605 ;
        RECT 553.355 3.915 553.685 4.245 ;
        RECT 553.355 2.555 553.685 2.885 ;
        RECT 553.355 1.195 553.685 1.525 ;
        RECT 553.355 -0.165 553.685 0.165 ;
        RECT 553.36 -8.32 553.68 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 554.715 10.715 555.045 11.045 ;
        RECT 554.715 9.355 555.045 9.685 ;
        RECT 554.715 7.995 555.045 8.325 ;
        RECT 554.715 6.635 555.045 6.965 ;
        RECT 554.715 5.275 555.045 5.605 ;
        RECT 554.715 3.915 555.045 4.245 ;
        RECT 554.715 2.555 555.045 2.885 ;
        RECT 554.715 1.195 555.045 1.525 ;
        RECT 554.715 -0.165 555.045 0.165 ;
        RECT 554.72 -8.32 555.04 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 556.075 10.715 556.405 11.045 ;
        RECT 556.075 9.355 556.405 9.685 ;
        RECT 556.075 7.995 556.405 8.325 ;
        RECT 556.075 6.635 556.405 6.965 ;
        RECT 556.075 5.275 556.405 5.605 ;
        RECT 556.075 3.915 556.405 4.245 ;
        RECT 556.075 2.555 556.405 2.885 ;
        RECT 556.075 1.195 556.405 1.525 ;
        RECT 556.075 -0.165 556.405 0.165 ;
        RECT 556.08 -8.32 556.4 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 557.435 10.715 557.765 11.045 ;
        RECT 557.435 9.355 557.765 9.685 ;
        RECT 557.435 7.995 557.765 8.325 ;
        RECT 557.435 6.635 557.765 6.965 ;
        RECT 557.435 5.275 557.765 5.605 ;
        RECT 557.435 3.915 557.765 4.245 ;
        RECT 557.435 2.555 557.765 2.885 ;
        RECT 557.435 1.195 557.765 1.525 ;
        RECT 557.435 -0.165 557.765 0.165 ;
        RECT 557.44 -8.32 557.76 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 558.795 10.715 559.125 11.045 ;
        RECT 558.795 9.355 559.125 9.685 ;
        RECT 558.795 7.995 559.125 8.325 ;
        RECT 558.795 6.635 559.125 6.965 ;
        RECT 558.795 5.275 559.125 5.605 ;
        RECT 558.795 3.915 559.125 4.245 ;
        RECT 558.795 2.555 559.125 2.885 ;
        RECT 558.795 1.195 559.125 1.525 ;
        RECT 558.795 -0.165 559.125 0.165 ;
        RECT 558.8 -8.32 559.12 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 560.155 10.715 560.485 11.045 ;
        RECT 560.155 9.355 560.485 9.685 ;
        RECT 560.155 7.995 560.485 8.325 ;
        RECT 560.155 6.635 560.485 6.965 ;
        RECT 560.155 5.275 560.485 5.605 ;
        RECT 560.155 3.915 560.485 4.245 ;
        RECT 560.155 2.555 560.485 2.885 ;
        RECT 560.155 1.195 560.485 1.525 ;
        RECT 560.155 -0.165 560.485 0.165 ;
        RECT 560.16 -8.32 560.48 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 561.515 10.715 561.845 11.045 ;
        RECT 561.515 9.355 561.845 9.685 ;
        RECT 561.515 7.995 561.845 8.325 ;
        RECT 561.515 6.635 561.845 6.965 ;
        RECT 561.515 5.275 561.845 5.605 ;
        RECT 561.515 3.915 561.845 4.245 ;
        RECT 561.515 2.555 561.845 2.885 ;
        RECT 561.515 1.195 561.845 1.525 ;
        RECT 561.515 -0.165 561.845 0.165 ;
        RECT 561.52 -8.32 561.84 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 562.875 10.715 563.205 11.045 ;
        RECT 562.875 9.355 563.205 9.685 ;
        RECT 562.875 7.995 563.205 8.325 ;
        RECT 562.875 6.635 563.205 6.965 ;
        RECT 562.875 5.275 563.205 5.605 ;
        RECT 562.875 3.915 563.205 4.245 ;
        RECT 562.875 2.555 563.205 2.885 ;
        RECT 562.875 1.195 563.205 1.525 ;
        RECT 562.875 -0.165 563.205 0.165 ;
        RECT 562.88 -8.32 563.2 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 564.235 10.715 564.565 11.045 ;
        RECT 564.235 9.355 564.565 9.685 ;
        RECT 564.235 7.995 564.565 8.325 ;
        RECT 564.235 6.635 564.565 6.965 ;
        RECT 564.235 5.275 564.565 5.605 ;
        RECT 564.235 3.915 564.565 4.245 ;
        RECT 564.235 2.555 564.565 2.885 ;
        RECT 564.235 1.195 564.565 1.525 ;
        RECT 564.235 -0.165 564.565 0.165 ;
        RECT 564.24 -8.32 564.56 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 565.595 10.715 565.925 11.045 ;
        RECT 565.595 9.355 565.925 9.685 ;
        RECT 565.595 7.995 565.925 8.325 ;
        RECT 565.595 6.635 565.925 6.965 ;
        RECT 565.595 5.275 565.925 5.605 ;
        RECT 565.595 3.915 565.925 4.245 ;
        RECT 565.595 2.555 565.925 2.885 ;
        RECT 565.595 1.195 565.925 1.525 ;
        RECT 565.595 -0.165 565.925 0.165 ;
        RECT 565.6 -8.32 565.92 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 566.955 10.715 567.285 11.045 ;
        RECT 566.955 9.355 567.285 9.685 ;
        RECT 566.955 7.995 567.285 8.325 ;
        RECT 566.955 6.635 567.285 6.965 ;
        RECT 566.955 5.275 567.285 5.605 ;
        RECT 566.955 3.915 567.285 4.245 ;
        RECT 566.955 2.555 567.285 2.885 ;
        RECT 566.955 1.195 567.285 1.525 ;
        RECT 566.955 -0.165 567.285 0.165 ;
        RECT 566.96 -8.32 567.28 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 568.315 10.715 568.645 11.045 ;
        RECT 568.315 9.355 568.645 9.685 ;
        RECT 568.315 7.995 568.645 8.325 ;
        RECT 568.315 6.635 568.645 6.965 ;
        RECT 568.315 5.275 568.645 5.605 ;
        RECT 568.315 3.915 568.645 4.245 ;
        RECT 568.315 2.555 568.645 2.885 ;
        RECT 568.315 1.195 568.645 1.525 ;
        RECT 568.315 -0.165 568.645 0.165 ;
        RECT 568.32 -8.32 568.64 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 569.675 10.715 570.005 11.045 ;
        RECT 569.675 9.355 570.005 9.685 ;
        RECT 569.675 7.995 570.005 8.325 ;
        RECT 569.675 6.635 570.005 6.965 ;
        RECT 569.675 5.275 570.005 5.605 ;
        RECT 569.675 3.915 570.005 4.245 ;
        RECT 569.675 2.555 570.005 2.885 ;
        RECT 569.675 1.195 570.005 1.525 ;
        RECT 569.675 -0.165 570.005 0.165 ;
        RECT 569.68 -8.32 570 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 571.035 10.715 571.365 11.045 ;
        RECT 571.035 9.355 571.365 9.685 ;
        RECT 571.035 7.995 571.365 8.325 ;
        RECT 571.035 6.635 571.365 6.965 ;
        RECT 571.035 5.275 571.365 5.605 ;
        RECT 571.035 3.915 571.365 4.245 ;
        RECT 571.035 2.555 571.365 2.885 ;
        RECT 571.035 1.195 571.365 1.525 ;
        RECT 571.035 -0.165 571.365 0.165 ;
        RECT 571.04 -8.32 571.36 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 572.395 10.715 572.725 11.045 ;
        RECT 572.395 9.355 572.725 9.685 ;
        RECT 572.395 7.995 572.725 8.325 ;
        RECT 572.395 6.635 572.725 6.965 ;
        RECT 572.395 5.275 572.725 5.605 ;
        RECT 572.395 3.915 572.725 4.245 ;
        RECT 572.395 2.555 572.725 2.885 ;
        RECT 572.395 1.195 572.725 1.525 ;
        RECT 572.395 -0.165 572.725 0.165 ;
        RECT 572.4 -8.32 572.72 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 573.755 10.715 574.085 11.045 ;
        RECT 573.755 9.355 574.085 9.685 ;
        RECT 573.755 7.995 574.085 8.325 ;
        RECT 573.755 6.635 574.085 6.965 ;
        RECT 573.755 5.275 574.085 5.605 ;
        RECT 573.755 3.915 574.085 4.245 ;
        RECT 573.755 2.555 574.085 2.885 ;
        RECT 573.755 1.195 574.085 1.525 ;
        RECT 573.755 -0.165 574.085 0.165 ;
        RECT 573.76 -8.32 574.08 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 575.115 10.715 575.445 11.045 ;
        RECT 575.115 9.355 575.445 9.685 ;
        RECT 575.115 7.995 575.445 8.325 ;
        RECT 575.115 6.635 575.445 6.965 ;
        RECT 575.115 5.275 575.445 5.605 ;
        RECT 575.115 3.915 575.445 4.245 ;
        RECT 575.115 2.555 575.445 2.885 ;
        RECT 575.115 1.195 575.445 1.525 ;
        RECT 575.115 -0.165 575.445 0.165 ;
        RECT 575.12 -8.32 575.44 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 576.475 10.715 576.805 11.045 ;
        RECT 576.475 9.355 576.805 9.685 ;
        RECT 576.475 7.995 576.805 8.325 ;
        RECT 576.475 6.635 576.805 6.965 ;
        RECT 576.475 5.275 576.805 5.605 ;
        RECT 576.475 3.915 576.805 4.245 ;
        RECT 576.475 2.555 576.805 2.885 ;
        RECT 576.475 1.195 576.805 1.525 ;
        RECT 576.475 -0.165 576.805 0.165 ;
        RECT 576.48 -8.32 576.8 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 577.835 10.715 578.165 11.045 ;
        RECT 577.835 9.355 578.165 9.685 ;
        RECT 577.835 7.995 578.165 8.325 ;
        RECT 577.835 6.635 578.165 6.965 ;
        RECT 577.835 5.275 578.165 5.605 ;
        RECT 577.835 3.915 578.165 4.245 ;
        RECT 577.835 2.555 578.165 2.885 ;
        RECT 577.835 1.195 578.165 1.525 ;
        RECT 577.835 -0.165 578.165 0.165 ;
        RECT 577.84 -8.32 578.16 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 579.195 10.715 579.525 11.045 ;
        RECT 579.195 9.355 579.525 9.685 ;
        RECT 579.195 7.995 579.525 8.325 ;
        RECT 579.195 6.635 579.525 6.965 ;
        RECT 579.195 5.275 579.525 5.605 ;
        RECT 579.195 3.915 579.525 4.245 ;
        RECT 579.195 2.555 579.525 2.885 ;
        RECT 579.195 1.195 579.525 1.525 ;
        RECT 579.195 -0.165 579.525 0.165 ;
        RECT 579.2 -8.32 579.52 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 580.555 10.715 580.885 11.045 ;
        RECT 580.555 9.355 580.885 9.685 ;
        RECT 580.555 7.995 580.885 8.325 ;
        RECT 580.555 6.635 580.885 6.965 ;
        RECT 580.555 5.275 580.885 5.605 ;
        RECT 580.555 3.915 580.885 4.245 ;
        RECT 580.555 2.555 580.885 2.885 ;
        RECT 580.555 1.195 580.885 1.525 ;
        RECT 580.555 -0.165 580.885 0.165 ;
        RECT 580.56 -8.32 580.88 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 581.915 10.715 582.245 11.045 ;
        RECT 581.915 9.355 582.245 9.685 ;
        RECT 581.915 7.995 582.245 8.325 ;
        RECT 581.915 6.635 582.245 6.965 ;
        RECT 581.915 5.275 582.245 5.605 ;
        RECT 581.915 3.915 582.245 4.245 ;
        RECT 581.915 2.555 582.245 2.885 ;
        RECT 581.915 1.195 582.245 1.525 ;
        RECT 581.915 -0.165 582.245 0.165 ;
        RECT 581.92 -8.32 582.24 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 583.275 10.715 583.605 11.045 ;
        RECT 583.275 9.355 583.605 9.685 ;
        RECT 583.275 7.995 583.605 8.325 ;
        RECT 583.275 6.635 583.605 6.965 ;
        RECT 583.275 5.275 583.605 5.605 ;
        RECT 583.275 3.915 583.605 4.245 ;
        RECT 583.275 2.555 583.605 2.885 ;
        RECT 583.275 1.195 583.605 1.525 ;
        RECT 583.275 -0.165 583.605 0.165 ;
        RECT 583.28 -8.32 583.6 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 584.635 10.715 584.965 11.045 ;
        RECT 584.635 9.355 584.965 9.685 ;
        RECT 584.635 7.995 584.965 8.325 ;
        RECT 584.635 6.635 584.965 6.965 ;
        RECT 584.635 5.275 584.965 5.605 ;
        RECT 584.635 3.915 584.965 4.245 ;
        RECT 584.635 2.555 584.965 2.885 ;
        RECT 584.635 1.195 584.965 1.525 ;
        RECT 584.635 -0.165 584.965 0.165 ;
        RECT 584.64 -8.32 584.96 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 585.995 10.715 586.325 11.045 ;
        RECT 585.995 9.355 586.325 9.685 ;
        RECT 585.995 7.995 586.325 8.325 ;
        RECT 585.995 6.635 586.325 6.965 ;
        RECT 585.995 5.275 586.325 5.605 ;
        RECT 585.995 3.915 586.325 4.245 ;
        RECT 585.995 2.555 586.325 2.885 ;
        RECT 585.995 1.195 586.325 1.525 ;
        RECT 585.995 -0.165 586.325 0.165 ;
        RECT 586 -8.32 586.32 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 587.355 10.715 587.685 11.045 ;
        RECT 587.355 9.355 587.685 9.685 ;
        RECT 587.355 7.995 587.685 8.325 ;
        RECT 587.355 6.635 587.685 6.965 ;
        RECT 587.355 5.275 587.685 5.605 ;
        RECT 587.355 3.915 587.685 4.245 ;
        RECT 587.355 2.555 587.685 2.885 ;
        RECT 587.355 1.195 587.685 1.525 ;
        RECT 587.355 -0.165 587.685 0.165 ;
        RECT 587.36 -8.32 587.68 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 588.715 10.715 589.045 11.045 ;
        RECT 588.715 9.355 589.045 9.685 ;
        RECT 588.715 7.995 589.045 8.325 ;
        RECT 588.715 6.635 589.045 6.965 ;
        RECT 588.715 5.275 589.045 5.605 ;
        RECT 588.715 3.915 589.045 4.245 ;
        RECT 588.715 2.555 589.045 2.885 ;
        RECT 588.715 1.195 589.045 1.525 ;
        RECT 588.715 -0.165 589.045 0.165 ;
        RECT 588.72 -8.32 589.04 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 590.075 10.715 590.405 11.045 ;
        RECT 590.075 9.355 590.405 9.685 ;
        RECT 590.075 7.995 590.405 8.325 ;
        RECT 590.075 6.635 590.405 6.965 ;
        RECT 590.075 5.275 590.405 5.605 ;
        RECT 590.075 3.915 590.405 4.245 ;
        RECT 590.075 2.555 590.405 2.885 ;
        RECT 590.075 1.195 590.405 1.525 ;
        RECT 590.075 -0.165 590.405 0.165 ;
        RECT 590.08 -8.32 590.4 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 591.435 10.715 591.765 11.045 ;
        RECT 591.435 9.355 591.765 9.685 ;
        RECT 591.435 7.995 591.765 8.325 ;
        RECT 591.435 6.635 591.765 6.965 ;
        RECT 591.435 5.275 591.765 5.605 ;
        RECT 591.435 3.915 591.765 4.245 ;
        RECT 591.435 2.555 591.765 2.885 ;
        RECT 591.435 1.195 591.765 1.525 ;
        RECT 591.435 -0.165 591.765 0.165 ;
        RECT 591.44 -8.32 591.76 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 592.795 10.715 593.125 11.045 ;
        RECT 592.795 9.355 593.125 9.685 ;
        RECT 592.795 7.995 593.125 8.325 ;
        RECT 592.795 6.635 593.125 6.965 ;
        RECT 592.795 5.275 593.125 5.605 ;
        RECT 592.795 3.915 593.125 4.245 ;
        RECT 592.795 2.555 593.125 2.885 ;
        RECT 592.795 1.195 593.125 1.525 ;
        RECT 592.795 -0.165 593.125 0.165 ;
        RECT 592.8 -8.32 593.12 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 594.155 10.715 594.485 11.045 ;
        RECT 594.155 9.355 594.485 9.685 ;
        RECT 594.155 7.995 594.485 8.325 ;
        RECT 594.155 6.635 594.485 6.965 ;
        RECT 594.155 5.275 594.485 5.605 ;
        RECT 594.155 3.915 594.485 4.245 ;
        RECT 594.155 2.555 594.485 2.885 ;
        RECT 594.155 1.195 594.485 1.525 ;
        RECT 594.155 -0.165 594.485 0.165 ;
        RECT 594.16 -8.32 594.48 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 595.515 10.715 595.845 11.045 ;
        RECT 595.515 9.355 595.845 9.685 ;
        RECT 595.515 7.995 595.845 8.325 ;
        RECT 595.515 6.635 595.845 6.965 ;
        RECT 595.515 5.275 595.845 5.605 ;
        RECT 595.515 3.915 595.845 4.245 ;
        RECT 595.515 2.555 595.845 2.885 ;
        RECT 595.515 1.195 595.845 1.525 ;
        RECT 595.515 -0.165 595.845 0.165 ;
        RECT 595.52 -8.32 595.84 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 596.875 10.715 597.205 11.045 ;
        RECT 596.875 9.355 597.205 9.685 ;
        RECT 596.875 7.995 597.205 8.325 ;
        RECT 596.875 6.635 597.205 6.965 ;
        RECT 596.875 5.275 597.205 5.605 ;
        RECT 596.875 3.915 597.205 4.245 ;
        RECT 596.875 2.555 597.205 2.885 ;
        RECT 596.875 1.195 597.205 1.525 ;
        RECT 596.875 -0.165 597.205 0.165 ;
        RECT 596.88 -8.32 597.2 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 598.235 10.715 598.565 11.045 ;
        RECT 598.235 9.355 598.565 9.685 ;
        RECT 598.235 7.995 598.565 8.325 ;
        RECT 598.235 6.635 598.565 6.965 ;
        RECT 598.235 5.275 598.565 5.605 ;
        RECT 598.235 3.915 598.565 4.245 ;
        RECT 598.235 2.555 598.565 2.885 ;
        RECT 598.235 1.195 598.565 1.525 ;
        RECT 598.235 -0.165 598.565 0.165 ;
        RECT 598.24 -8.32 598.56 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 599.595 10.715 599.925 11.045 ;
        RECT 599.595 9.355 599.925 9.685 ;
        RECT 599.595 7.995 599.925 8.325 ;
        RECT 599.595 6.635 599.925 6.965 ;
        RECT 599.595 5.275 599.925 5.605 ;
        RECT 599.595 3.915 599.925 4.245 ;
        RECT 599.595 2.555 599.925 2.885 ;
        RECT 599.595 1.195 599.925 1.525 ;
        RECT 599.595 -0.165 599.925 0.165 ;
        RECT 599.6 -8.32 599.92 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 600.955 10.715 601.285 11.045 ;
        RECT 600.955 9.355 601.285 9.685 ;
        RECT 600.955 7.995 601.285 8.325 ;
        RECT 600.955 6.635 601.285 6.965 ;
        RECT 600.955 5.275 601.285 5.605 ;
        RECT 600.955 3.915 601.285 4.245 ;
        RECT 600.955 2.555 601.285 2.885 ;
        RECT 600.955 1.195 601.285 1.525 ;
        RECT 600.955 -0.165 601.285 0.165 ;
        RECT 600.96 -8.32 601.28 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 602.315 10.715 602.645 11.045 ;
        RECT 602.315 9.355 602.645 9.685 ;
        RECT 602.315 7.995 602.645 8.325 ;
        RECT 602.315 6.635 602.645 6.965 ;
        RECT 602.315 5.275 602.645 5.605 ;
        RECT 602.315 3.915 602.645 4.245 ;
        RECT 602.315 2.555 602.645 2.885 ;
        RECT 602.315 1.195 602.645 1.525 ;
        RECT 602.315 -0.165 602.645 0.165 ;
        RECT 602.32 -8.32 602.64 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 603.675 10.715 604.005 11.045 ;
        RECT 603.675 9.355 604.005 9.685 ;
        RECT 603.675 7.995 604.005 8.325 ;
        RECT 603.675 6.635 604.005 6.965 ;
        RECT 603.675 5.275 604.005 5.605 ;
        RECT 603.675 3.915 604.005 4.245 ;
        RECT 603.675 2.555 604.005 2.885 ;
        RECT 603.675 1.195 604.005 1.525 ;
        RECT 603.675 -0.165 604.005 0.165 ;
        RECT 603.68 -8.32 604 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 605.035 10.715 605.365 11.045 ;
        RECT 605.035 9.355 605.365 9.685 ;
        RECT 605.035 7.995 605.365 8.325 ;
        RECT 605.035 6.635 605.365 6.965 ;
        RECT 605.035 5.275 605.365 5.605 ;
        RECT 605.035 3.915 605.365 4.245 ;
        RECT 605.035 2.555 605.365 2.885 ;
        RECT 605.035 1.195 605.365 1.525 ;
        RECT 605.035 -0.165 605.365 0.165 ;
        RECT 605.04 -8.32 605.36 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 606.395 10.715 606.725 11.045 ;
        RECT 606.395 9.355 606.725 9.685 ;
        RECT 606.395 7.995 606.725 8.325 ;
        RECT 606.395 6.635 606.725 6.965 ;
        RECT 606.395 5.275 606.725 5.605 ;
        RECT 606.395 3.915 606.725 4.245 ;
        RECT 606.395 2.555 606.725 2.885 ;
        RECT 606.395 1.195 606.725 1.525 ;
        RECT 606.395 -0.165 606.725 0.165 ;
        RECT 606.4 -8.32 606.72 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 607.755 10.715 608.085 11.045 ;
        RECT 607.755 9.355 608.085 9.685 ;
        RECT 607.755 7.995 608.085 8.325 ;
        RECT 607.755 6.635 608.085 6.965 ;
        RECT 607.755 5.275 608.085 5.605 ;
        RECT 607.755 3.915 608.085 4.245 ;
        RECT 607.755 2.555 608.085 2.885 ;
        RECT 607.755 1.195 608.085 1.525 ;
        RECT 607.755 -0.165 608.085 0.165 ;
        RECT 607.76 -8.32 608.08 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 609.115 10.715 609.445 11.045 ;
        RECT 609.115 9.355 609.445 9.685 ;
        RECT 609.115 7.995 609.445 8.325 ;
        RECT 609.115 6.635 609.445 6.965 ;
        RECT 609.115 5.275 609.445 5.605 ;
        RECT 609.115 3.915 609.445 4.245 ;
        RECT 609.115 2.555 609.445 2.885 ;
        RECT 609.115 1.195 609.445 1.525 ;
        RECT 609.115 -0.165 609.445 0.165 ;
        RECT 609.12 -8.32 609.44 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 610.475 10.715 610.805 11.045 ;
        RECT 610.475 9.355 610.805 9.685 ;
        RECT 610.475 7.995 610.805 8.325 ;
        RECT 610.475 6.635 610.805 6.965 ;
        RECT 610.475 5.275 610.805 5.605 ;
        RECT 610.475 3.915 610.805 4.245 ;
        RECT 610.475 2.555 610.805 2.885 ;
        RECT 610.475 1.195 610.805 1.525 ;
        RECT 610.475 -0.165 610.805 0.165 ;
        RECT 610.48 -8.32 610.8 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 611.835 10.715 612.165 11.045 ;
        RECT 611.835 9.355 612.165 9.685 ;
        RECT 611.835 7.995 612.165 8.325 ;
        RECT 611.835 6.635 612.165 6.965 ;
        RECT 611.835 5.275 612.165 5.605 ;
        RECT 611.835 3.915 612.165 4.245 ;
        RECT 611.835 2.555 612.165 2.885 ;
        RECT 611.835 1.195 612.165 1.525 ;
        RECT 611.835 -0.165 612.165 0.165 ;
        RECT 611.84 -8.32 612.16 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 613.195 10.715 613.525 11.045 ;
        RECT 613.195 9.355 613.525 9.685 ;
        RECT 613.195 7.995 613.525 8.325 ;
        RECT 613.195 6.635 613.525 6.965 ;
        RECT 613.195 5.275 613.525 5.605 ;
        RECT 613.195 3.915 613.525 4.245 ;
        RECT 613.195 2.555 613.525 2.885 ;
        RECT 613.195 1.195 613.525 1.525 ;
        RECT 613.195 -0.165 613.525 0.165 ;
        RECT 613.2 -8.32 613.52 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 614.555 10.715 614.885 11.045 ;
        RECT 614.555 9.355 614.885 9.685 ;
        RECT 614.555 7.995 614.885 8.325 ;
        RECT 614.555 6.635 614.885 6.965 ;
        RECT 614.555 5.275 614.885 5.605 ;
        RECT 614.555 3.915 614.885 4.245 ;
        RECT 614.555 2.555 614.885 2.885 ;
        RECT 614.555 1.195 614.885 1.525 ;
        RECT 614.555 -0.165 614.885 0.165 ;
        RECT 614.56 -8.32 614.88 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 615.915 10.715 616.245 11.045 ;
        RECT 615.915 9.355 616.245 9.685 ;
        RECT 615.915 7.995 616.245 8.325 ;
        RECT 615.915 6.635 616.245 6.965 ;
        RECT 615.915 5.275 616.245 5.605 ;
        RECT 615.915 3.915 616.245 4.245 ;
        RECT 615.915 2.555 616.245 2.885 ;
        RECT 615.915 1.195 616.245 1.525 ;
        RECT 615.915 -0.165 616.245 0.165 ;
        RECT 615.92 -8.32 616.24 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 617.275 10.715 617.605 11.045 ;
        RECT 617.275 9.355 617.605 9.685 ;
        RECT 617.275 7.995 617.605 8.325 ;
        RECT 617.275 6.635 617.605 6.965 ;
        RECT 617.275 5.275 617.605 5.605 ;
        RECT 617.275 3.915 617.605 4.245 ;
        RECT 617.275 2.555 617.605 2.885 ;
        RECT 617.275 1.195 617.605 1.525 ;
        RECT 617.275 -0.165 617.605 0.165 ;
        RECT 617.28 -8.32 617.6 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 618.635 10.715 618.965 11.045 ;
        RECT 618.635 9.355 618.965 9.685 ;
        RECT 618.635 7.995 618.965 8.325 ;
        RECT 618.635 6.635 618.965 6.965 ;
        RECT 618.635 5.275 618.965 5.605 ;
        RECT 618.635 3.915 618.965 4.245 ;
        RECT 618.635 2.555 618.965 2.885 ;
        RECT 618.635 1.195 618.965 1.525 ;
        RECT 618.635 -0.165 618.965 0.165 ;
        RECT 618.64 -8.32 618.96 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 619.995 10.715 620.325 11.045 ;
        RECT 619.995 9.355 620.325 9.685 ;
        RECT 619.995 7.995 620.325 8.325 ;
        RECT 619.995 6.635 620.325 6.965 ;
        RECT 619.995 5.275 620.325 5.605 ;
        RECT 619.995 3.915 620.325 4.245 ;
        RECT 619.995 2.555 620.325 2.885 ;
        RECT 619.995 1.195 620.325 1.525 ;
        RECT 619.995 -0.165 620.325 0.165 ;
        RECT 620 -8.32 620.32 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 621.355 10.715 621.685 11.045 ;
        RECT 621.355 9.355 621.685 9.685 ;
        RECT 621.355 7.995 621.685 8.325 ;
        RECT 621.355 6.635 621.685 6.965 ;
        RECT 621.355 5.275 621.685 5.605 ;
        RECT 621.355 3.915 621.685 4.245 ;
        RECT 621.355 2.555 621.685 2.885 ;
        RECT 621.355 1.195 621.685 1.525 ;
        RECT 621.355 -0.165 621.685 0.165 ;
        RECT 621.36 -8.32 621.68 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 622.715 10.715 623.045 11.045 ;
        RECT 622.715 9.355 623.045 9.685 ;
        RECT 622.715 7.995 623.045 8.325 ;
        RECT 622.715 6.635 623.045 6.965 ;
        RECT 622.715 5.275 623.045 5.605 ;
        RECT 622.715 3.915 623.045 4.245 ;
        RECT 622.715 2.555 623.045 2.885 ;
        RECT 622.715 1.195 623.045 1.525 ;
        RECT 622.715 -0.165 623.045 0.165 ;
        RECT 622.72 -8.32 623.04 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 624.075 10.715 624.405 11.045 ;
        RECT 624.075 9.355 624.405 9.685 ;
        RECT 624.075 7.995 624.405 8.325 ;
        RECT 624.075 6.635 624.405 6.965 ;
        RECT 624.075 5.275 624.405 5.605 ;
        RECT 624.075 3.915 624.405 4.245 ;
        RECT 624.075 2.555 624.405 2.885 ;
        RECT 624.075 1.195 624.405 1.525 ;
        RECT 624.075 -0.165 624.405 0.165 ;
        RECT 624.08 -8.32 624.4 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 625.435 10.715 625.765 11.045 ;
        RECT 625.435 9.355 625.765 9.685 ;
        RECT 625.435 7.995 625.765 8.325 ;
        RECT 625.435 6.635 625.765 6.965 ;
        RECT 625.435 5.275 625.765 5.605 ;
        RECT 625.435 3.915 625.765 4.245 ;
        RECT 625.435 2.555 625.765 2.885 ;
        RECT 625.435 1.195 625.765 1.525 ;
        RECT 625.435 -0.165 625.765 0.165 ;
        RECT 625.44 -8.32 625.76 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 626.795 10.715 627.125 11.045 ;
        RECT 626.795 9.355 627.125 9.685 ;
        RECT 626.795 7.995 627.125 8.325 ;
        RECT 626.795 6.635 627.125 6.965 ;
        RECT 626.795 5.275 627.125 5.605 ;
        RECT 626.795 3.915 627.125 4.245 ;
        RECT 626.795 2.555 627.125 2.885 ;
        RECT 626.795 1.195 627.125 1.525 ;
        RECT 626.795 -0.165 627.125 0.165 ;
        RECT 626.8 -8.32 627.12 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 628.155 10.715 628.485 11.045 ;
        RECT 628.155 9.355 628.485 9.685 ;
        RECT 628.155 7.995 628.485 8.325 ;
        RECT 628.155 6.635 628.485 6.965 ;
        RECT 628.155 5.275 628.485 5.605 ;
        RECT 628.155 3.915 628.485 4.245 ;
        RECT 628.155 2.555 628.485 2.885 ;
        RECT 628.155 1.195 628.485 1.525 ;
        RECT 628.155 -0.165 628.485 0.165 ;
        RECT 628.16 -8.32 628.48 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 629.515 10.715 629.845 11.045 ;
        RECT 629.515 9.355 629.845 9.685 ;
        RECT 629.515 7.995 629.845 8.325 ;
        RECT 629.515 6.635 629.845 6.965 ;
        RECT 629.515 5.275 629.845 5.605 ;
        RECT 629.515 3.915 629.845 4.245 ;
        RECT 629.515 2.555 629.845 2.885 ;
        RECT 629.515 1.195 629.845 1.525 ;
        RECT 629.515 -0.165 629.845 0.165 ;
        RECT 629.52 -8.32 629.84 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 630.875 10.715 631.205 11.045 ;
        RECT 630.875 9.355 631.205 9.685 ;
        RECT 630.875 7.995 631.205 8.325 ;
        RECT 630.875 6.635 631.205 6.965 ;
        RECT 630.875 5.275 631.205 5.605 ;
        RECT 630.875 3.915 631.205 4.245 ;
        RECT 630.875 2.555 631.205 2.885 ;
        RECT 630.875 1.195 631.205 1.525 ;
        RECT 630.875 -0.165 631.205 0.165 ;
        RECT 630.88 -8.32 631.2 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 632.235 10.715 632.565 11.045 ;
        RECT 632.235 9.355 632.565 9.685 ;
        RECT 632.235 7.995 632.565 8.325 ;
        RECT 632.235 6.635 632.565 6.965 ;
        RECT 632.235 5.275 632.565 5.605 ;
        RECT 632.235 3.915 632.565 4.245 ;
        RECT 632.235 2.555 632.565 2.885 ;
        RECT 632.235 1.195 632.565 1.525 ;
        RECT 632.235 -0.165 632.565 0.165 ;
        RECT 632.24 -8.32 632.56 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 633.595 9.355 633.925 9.685 ;
        RECT 633.595 7.995 633.925 8.325 ;
        RECT 633.595 6.635 633.925 6.965 ;
        RECT 633.595 5.275 633.925 5.605 ;
        RECT 633.595 3.915 633.925 4.245 ;
        RECT 633.595 2.555 633.925 2.885 ;
        RECT 633.595 1.195 633.925 1.525 ;
        RECT 633.595 -0.165 633.925 0.165 ;
        RECT 633.6 -8.32 633.92 15.8 ;
        RECT 633.595 10.715 633.925 11.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 362.955 10.715 363.285 11.045 ;
        RECT 362.955 9.355 363.285 9.685 ;
        RECT 362.955 7.995 363.285 8.325 ;
        RECT 362.955 6.635 363.285 6.965 ;
        RECT 362.955 5.275 363.285 5.605 ;
        RECT 362.955 3.915 363.285 4.245 ;
        RECT 362.955 2.555 363.285 2.885 ;
        RECT 362.955 1.195 363.285 1.525 ;
        RECT 362.955 -0.165 363.285 0.165 ;
        RECT 362.96 -8.32 363.28 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 364.315 10.715 364.645 11.045 ;
        RECT 364.315 9.355 364.645 9.685 ;
        RECT 364.315 7.995 364.645 8.325 ;
        RECT 364.315 6.635 364.645 6.965 ;
        RECT 364.315 5.275 364.645 5.605 ;
        RECT 364.315 3.915 364.645 4.245 ;
        RECT 364.315 2.555 364.645 2.885 ;
        RECT 364.315 1.195 364.645 1.525 ;
        RECT 364.315 -0.165 364.645 0.165 ;
        RECT 364.32 -8.32 364.64 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 365.675 10.715 366.005 11.045 ;
        RECT 365.675 9.355 366.005 9.685 ;
        RECT 365.675 7.995 366.005 8.325 ;
        RECT 365.675 6.635 366.005 6.965 ;
        RECT 365.675 5.275 366.005 5.605 ;
        RECT 365.675 3.915 366.005 4.245 ;
        RECT 365.675 2.555 366.005 2.885 ;
        RECT 365.675 1.195 366.005 1.525 ;
        RECT 365.675 -0.165 366.005 0.165 ;
        RECT 365.68 -8.32 366 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 367.035 10.715 367.365 11.045 ;
        RECT 367.035 9.355 367.365 9.685 ;
        RECT 367.035 7.995 367.365 8.325 ;
        RECT 367.035 6.635 367.365 6.965 ;
        RECT 367.035 5.275 367.365 5.605 ;
        RECT 367.035 3.915 367.365 4.245 ;
        RECT 367.035 2.555 367.365 2.885 ;
        RECT 367.035 1.195 367.365 1.525 ;
        RECT 367.035 -0.165 367.365 0.165 ;
        RECT 367.04 -8.32 367.36 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 368.395 10.715 368.725 11.045 ;
        RECT 368.395 9.355 368.725 9.685 ;
        RECT 368.395 7.995 368.725 8.325 ;
        RECT 368.395 6.635 368.725 6.965 ;
        RECT 368.395 5.275 368.725 5.605 ;
        RECT 368.395 3.915 368.725 4.245 ;
        RECT 368.395 2.555 368.725 2.885 ;
        RECT 368.395 1.195 368.725 1.525 ;
        RECT 368.395 -0.165 368.725 0.165 ;
        RECT 368.4 -8.32 368.72 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 369.755 10.715 370.085 11.045 ;
        RECT 369.755 9.355 370.085 9.685 ;
        RECT 369.755 7.995 370.085 8.325 ;
        RECT 369.755 6.635 370.085 6.965 ;
        RECT 369.755 5.275 370.085 5.605 ;
        RECT 369.755 3.915 370.085 4.245 ;
        RECT 369.755 2.555 370.085 2.885 ;
        RECT 369.755 1.195 370.085 1.525 ;
        RECT 369.755 -0.165 370.085 0.165 ;
        RECT 369.76 -8.32 370.08 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 371.115 10.715 371.445 11.045 ;
        RECT 371.115 9.355 371.445 9.685 ;
        RECT 371.115 7.995 371.445 8.325 ;
        RECT 371.115 6.635 371.445 6.965 ;
        RECT 371.115 5.275 371.445 5.605 ;
        RECT 371.115 3.915 371.445 4.245 ;
        RECT 371.115 2.555 371.445 2.885 ;
        RECT 371.115 1.195 371.445 1.525 ;
        RECT 371.115 -0.165 371.445 0.165 ;
        RECT 371.12 -8.32 371.44 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 372.475 10.715 372.805 11.045 ;
        RECT 372.475 9.355 372.805 9.685 ;
        RECT 372.475 7.995 372.805 8.325 ;
        RECT 372.475 6.635 372.805 6.965 ;
        RECT 372.475 5.275 372.805 5.605 ;
        RECT 372.475 3.915 372.805 4.245 ;
        RECT 372.475 2.555 372.805 2.885 ;
        RECT 372.475 1.195 372.805 1.525 ;
        RECT 372.475 -0.165 372.805 0.165 ;
        RECT 372.48 -8.32 372.8 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 373.835 10.715 374.165 11.045 ;
        RECT 373.835 9.355 374.165 9.685 ;
        RECT 373.835 7.995 374.165 8.325 ;
        RECT 373.835 6.635 374.165 6.965 ;
        RECT 373.835 5.275 374.165 5.605 ;
        RECT 373.835 3.915 374.165 4.245 ;
        RECT 373.835 2.555 374.165 2.885 ;
        RECT 373.835 1.195 374.165 1.525 ;
        RECT 373.835 -0.165 374.165 0.165 ;
        RECT 373.84 -8.32 374.16 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 375.195 10.715 375.525 11.045 ;
        RECT 375.195 9.355 375.525 9.685 ;
        RECT 375.195 7.995 375.525 8.325 ;
        RECT 375.195 6.635 375.525 6.965 ;
        RECT 375.195 5.275 375.525 5.605 ;
        RECT 375.195 3.915 375.525 4.245 ;
        RECT 375.195 2.555 375.525 2.885 ;
        RECT 375.195 1.195 375.525 1.525 ;
        RECT 375.195 -0.165 375.525 0.165 ;
        RECT 375.2 -8.32 375.52 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 376.555 10.715 376.885 11.045 ;
        RECT 376.555 9.355 376.885 9.685 ;
        RECT 376.555 7.995 376.885 8.325 ;
        RECT 376.555 6.635 376.885 6.965 ;
        RECT 376.555 5.275 376.885 5.605 ;
        RECT 376.555 3.915 376.885 4.245 ;
        RECT 376.555 2.555 376.885 2.885 ;
        RECT 376.555 1.195 376.885 1.525 ;
        RECT 376.555 -0.165 376.885 0.165 ;
        RECT 376.56 -8.32 376.88 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 377.915 10.715 378.245 11.045 ;
        RECT 377.915 9.355 378.245 9.685 ;
        RECT 377.915 7.995 378.245 8.325 ;
        RECT 377.915 6.635 378.245 6.965 ;
        RECT 377.915 5.275 378.245 5.605 ;
        RECT 377.915 3.915 378.245 4.245 ;
        RECT 377.915 2.555 378.245 2.885 ;
        RECT 377.915 1.195 378.245 1.525 ;
        RECT 377.915 -0.165 378.245 0.165 ;
        RECT 377.92 -8.32 378.24 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 379.275 10.715 379.605 11.045 ;
        RECT 379.275 9.355 379.605 9.685 ;
        RECT 379.275 7.995 379.605 8.325 ;
        RECT 379.275 6.635 379.605 6.965 ;
        RECT 379.275 5.275 379.605 5.605 ;
        RECT 379.275 3.915 379.605 4.245 ;
        RECT 379.275 2.555 379.605 2.885 ;
        RECT 379.275 1.195 379.605 1.525 ;
        RECT 379.275 -0.165 379.605 0.165 ;
        RECT 379.28 -8.32 379.6 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 380.635 10.715 380.965 11.045 ;
        RECT 380.635 9.355 380.965 9.685 ;
        RECT 380.635 7.995 380.965 8.325 ;
        RECT 380.635 6.635 380.965 6.965 ;
        RECT 380.635 5.275 380.965 5.605 ;
        RECT 380.635 3.915 380.965 4.245 ;
        RECT 380.635 2.555 380.965 2.885 ;
        RECT 380.635 1.195 380.965 1.525 ;
        RECT 380.635 -0.165 380.965 0.165 ;
        RECT 380.64 -8.32 380.96 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 381.995 10.715 382.325 11.045 ;
        RECT 381.995 9.355 382.325 9.685 ;
        RECT 381.995 7.995 382.325 8.325 ;
        RECT 381.995 6.635 382.325 6.965 ;
        RECT 381.995 5.275 382.325 5.605 ;
        RECT 381.995 3.915 382.325 4.245 ;
        RECT 381.995 2.555 382.325 2.885 ;
        RECT 381.995 1.195 382.325 1.525 ;
        RECT 381.995 -0.165 382.325 0.165 ;
        RECT 382 -8.32 382.32 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 383.355 10.715 383.685 11.045 ;
        RECT 383.355 9.355 383.685 9.685 ;
        RECT 383.355 7.995 383.685 8.325 ;
        RECT 383.355 6.635 383.685 6.965 ;
        RECT 383.355 5.275 383.685 5.605 ;
        RECT 383.355 3.915 383.685 4.245 ;
        RECT 383.355 2.555 383.685 2.885 ;
        RECT 383.355 1.195 383.685 1.525 ;
        RECT 383.355 -0.165 383.685 0.165 ;
        RECT 383.36 -8.32 383.68 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 384.715 10.715 385.045 11.045 ;
        RECT 384.715 9.355 385.045 9.685 ;
        RECT 384.715 7.995 385.045 8.325 ;
        RECT 384.715 6.635 385.045 6.965 ;
        RECT 384.715 5.275 385.045 5.605 ;
        RECT 384.715 3.915 385.045 4.245 ;
        RECT 384.715 2.555 385.045 2.885 ;
        RECT 384.715 1.195 385.045 1.525 ;
        RECT 384.715 -0.165 385.045 0.165 ;
        RECT 384.72 -8.32 385.04 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 386.075 10.715 386.405 11.045 ;
        RECT 386.075 9.355 386.405 9.685 ;
        RECT 386.075 7.995 386.405 8.325 ;
        RECT 386.075 6.635 386.405 6.965 ;
        RECT 386.075 5.275 386.405 5.605 ;
        RECT 386.075 3.915 386.405 4.245 ;
        RECT 386.075 2.555 386.405 2.885 ;
        RECT 386.075 1.195 386.405 1.525 ;
        RECT 386.075 -0.165 386.405 0.165 ;
        RECT 386.08 -8.32 386.4 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 387.435 10.715 387.765 11.045 ;
        RECT 387.435 9.355 387.765 9.685 ;
        RECT 387.435 7.995 387.765 8.325 ;
        RECT 387.435 6.635 387.765 6.965 ;
        RECT 387.435 5.275 387.765 5.605 ;
        RECT 387.435 3.915 387.765 4.245 ;
        RECT 387.435 2.555 387.765 2.885 ;
        RECT 387.435 1.195 387.765 1.525 ;
        RECT 387.435 -0.165 387.765 0.165 ;
        RECT 387.44 -8.32 387.76 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 388.795 10.715 389.125 11.045 ;
        RECT 388.795 9.355 389.125 9.685 ;
        RECT 388.795 7.995 389.125 8.325 ;
        RECT 388.795 6.635 389.125 6.965 ;
        RECT 388.795 5.275 389.125 5.605 ;
        RECT 388.795 3.915 389.125 4.245 ;
        RECT 388.795 2.555 389.125 2.885 ;
        RECT 388.795 1.195 389.125 1.525 ;
        RECT 388.795 -0.165 389.125 0.165 ;
        RECT 388.8 -8.32 389.12 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 390.155 10.715 390.485 11.045 ;
        RECT 390.155 9.355 390.485 9.685 ;
        RECT 390.155 7.995 390.485 8.325 ;
        RECT 390.155 6.635 390.485 6.965 ;
        RECT 390.155 5.275 390.485 5.605 ;
        RECT 390.155 3.915 390.485 4.245 ;
        RECT 390.155 2.555 390.485 2.885 ;
        RECT 390.155 1.195 390.485 1.525 ;
        RECT 390.155 -0.165 390.485 0.165 ;
        RECT 390.16 -8.32 390.48 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 391.515 10.715 391.845 11.045 ;
        RECT 391.515 9.355 391.845 9.685 ;
        RECT 391.515 7.995 391.845 8.325 ;
        RECT 391.515 6.635 391.845 6.965 ;
        RECT 391.515 5.275 391.845 5.605 ;
        RECT 391.515 3.915 391.845 4.245 ;
        RECT 391.515 2.555 391.845 2.885 ;
        RECT 391.515 1.195 391.845 1.525 ;
        RECT 391.515 -0.165 391.845 0.165 ;
        RECT 391.52 -8.32 391.84 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 392.875 10.715 393.205 11.045 ;
        RECT 392.875 9.355 393.205 9.685 ;
        RECT 392.875 7.995 393.205 8.325 ;
        RECT 392.875 6.635 393.205 6.965 ;
        RECT 392.875 5.275 393.205 5.605 ;
        RECT 392.875 3.915 393.205 4.245 ;
        RECT 392.875 2.555 393.205 2.885 ;
        RECT 392.875 1.195 393.205 1.525 ;
        RECT 392.875 -0.165 393.205 0.165 ;
        RECT 392.88 -8.32 393.2 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 394.235 10.715 394.565 11.045 ;
        RECT 394.235 9.355 394.565 9.685 ;
        RECT 394.235 7.995 394.565 8.325 ;
        RECT 394.235 6.635 394.565 6.965 ;
        RECT 394.235 5.275 394.565 5.605 ;
        RECT 394.235 3.915 394.565 4.245 ;
        RECT 394.235 2.555 394.565 2.885 ;
        RECT 394.235 1.195 394.565 1.525 ;
        RECT 394.235 -0.165 394.565 0.165 ;
        RECT 394.24 -8.32 394.56 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 395.595 10.715 395.925 11.045 ;
        RECT 395.595 9.355 395.925 9.685 ;
        RECT 395.595 7.995 395.925 8.325 ;
        RECT 395.595 6.635 395.925 6.965 ;
        RECT 395.595 5.275 395.925 5.605 ;
        RECT 395.595 3.915 395.925 4.245 ;
        RECT 395.595 2.555 395.925 2.885 ;
        RECT 395.595 1.195 395.925 1.525 ;
        RECT 395.595 -0.165 395.925 0.165 ;
        RECT 395.6 -8.32 395.92 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 396.955 10.715 397.285 11.045 ;
        RECT 396.955 9.355 397.285 9.685 ;
        RECT 396.955 7.995 397.285 8.325 ;
        RECT 396.955 6.635 397.285 6.965 ;
        RECT 396.955 5.275 397.285 5.605 ;
        RECT 396.955 3.915 397.285 4.245 ;
        RECT 396.955 2.555 397.285 2.885 ;
        RECT 396.955 1.195 397.285 1.525 ;
        RECT 396.955 -0.165 397.285 0.165 ;
        RECT 396.96 -8.32 397.28 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 398.315 10.715 398.645 11.045 ;
        RECT 398.315 9.355 398.645 9.685 ;
        RECT 398.315 7.995 398.645 8.325 ;
        RECT 398.315 6.635 398.645 6.965 ;
        RECT 398.315 5.275 398.645 5.605 ;
        RECT 398.315 3.915 398.645 4.245 ;
        RECT 398.315 2.555 398.645 2.885 ;
        RECT 398.315 1.195 398.645 1.525 ;
        RECT 398.315 -0.165 398.645 0.165 ;
        RECT 398.32 -8.32 398.64 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 399.675 10.715 400.005 11.045 ;
        RECT 399.675 9.355 400.005 9.685 ;
        RECT 399.675 7.995 400.005 8.325 ;
        RECT 399.675 6.635 400.005 6.965 ;
        RECT 399.675 5.275 400.005 5.605 ;
        RECT 399.675 3.915 400.005 4.245 ;
        RECT 399.675 2.555 400.005 2.885 ;
        RECT 399.675 1.195 400.005 1.525 ;
        RECT 399.675 -0.165 400.005 0.165 ;
        RECT 399.68 -8.32 400 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 401.035 10.715 401.365 11.045 ;
        RECT 401.035 9.355 401.365 9.685 ;
        RECT 401.035 7.995 401.365 8.325 ;
        RECT 401.035 6.635 401.365 6.965 ;
        RECT 401.035 5.275 401.365 5.605 ;
        RECT 401.035 3.915 401.365 4.245 ;
        RECT 401.035 2.555 401.365 2.885 ;
        RECT 401.035 1.195 401.365 1.525 ;
        RECT 401.035 -0.165 401.365 0.165 ;
        RECT 401.04 -8.32 401.36 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 402.395 10.715 402.725 11.045 ;
        RECT 402.395 9.355 402.725 9.685 ;
        RECT 402.395 7.995 402.725 8.325 ;
        RECT 402.395 6.635 402.725 6.965 ;
        RECT 402.395 5.275 402.725 5.605 ;
        RECT 402.395 3.915 402.725 4.245 ;
        RECT 402.395 2.555 402.725 2.885 ;
        RECT 402.395 1.195 402.725 1.525 ;
        RECT 402.395 -0.165 402.725 0.165 ;
        RECT 402.4 -8.32 402.72 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 403.755 10.715 404.085 11.045 ;
        RECT 403.755 9.355 404.085 9.685 ;
        RECT 403.755 7.995 404.085 8.325 ;
        RECT 403.755 6.635 404.085 6.965 ;
        RECT 403.755 5.275 404.085 5.605 ;
        RECT 403.755 3.915 404.085 4.245 ;
        RECT 403.755 2.555 404.085 2.885 ;
        RECT 403.755 1.195 404.085 1.525 ;
        RECT 403.755 -0.165 404.085 0.165 ;
        RECT 403.76 -8.32 404.08 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 405.115 10.715 405.445 11.045 ;
        RECT 405.115 9.355 405.445 9.685 ;
        RECT 405.115 7.995 405.445 8.325 ;
        RECT 405.115 6.635 405.445 6.965 ;
        RECT 405.115 5.275 405.445 5.605 ;
        RECT 405.115 3.915 405.445 4.245 ;
        RECT 405.115 2.555 405.445 2.885 ;
        RECT 405.115 1.195 405.445 1.525 ;
        RECT 405.115 -0.165 405.445 0.165 ;
        RECT 405.12 -8.32 405.44 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 406.475 10.715 406.805 11.045 ;
        RECT 406.475 9.355 406.805 9.685 ;
        RECT 406.475 7.995 406.805 8.325 ;
        RECT 406.475 6.635 406.805 6.965 ;
        RECT 406.475 5.275 406.805 5.605 ;
        RECT 406.475 3.915 406.805 4.245 ;
        RECT 406.475 2.555 406.805 2.885 ;
        RECT 406.475 1.195 406.805 1.525 ;
        RECT 406.475 -0.165 406.805 0.165 ;
        RECT 406.48 -8.32 406.8 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 407.835 10.715 408.165 11.045 ;
        RECT 407.835 9.355 408.165 9.685 ;
        RECT 407.835 7.995 408.165 8.325 ;
        RECT 407.835 6.635 408.165 6.965 ;
        RECT 407.835 5.275 408.165 5.605 ;
        RECT 407.835 3.915 408.165 4.245 ;
        RECT 407.835 2.555 408.165 2.885 ;
        RECT 407.835 1.195 408.165 1.525 ;
        RECT 407.835 -0.165 408.165 0.165 ;
        RECT 407.84 -8.32 408.16 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 409.195 10.715 409.525 11.045 ;
        RECT 409.195 9.355 409.525 9.685 ;
        RECT 409.195 7.995 409.525 8.325 ;
        RECT 409.195 6.635 409.525 6.965 ;
        RECT 409.195 5.275 409.525 5.605 ;
        RECT 409.195 3.915 409.525 4.245 ;
        RECT 409.195 2.555 409.525 2.885 ;
        RECT 409.195 1.195 409.525 1.525 ;
        RECT 409.195 -0.165 409.525 0.165 ;
        RECT 409.2 -8.32 409.52 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 410.555 10.715 410.885 11.045 ;
        RECT 410.555 9.355 410.885 9.685 ;
        RECT 410.555 7.995 410.885 8.325 ;
        RECT 410.555 6.635 410.885 6.965 ;
        RECT 410.555 5.275 410.885 5.605 ;
        RECT 410.555 3.915 410.885 4.245 ;
        RECT 410.555 2.555 410.885 2.885 ;
        RECT 410.555 1.195 410.885 1.525 ;
        RECT 410.555 -0.165 410.885 0.165 ;
        RECT 410.56 -8.32 410.88 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 411.915 10.715 412.245 11.045 ;
        RECT 411.915 9.355 412.245 9.685 ;
        RECT 411.915 7.995 412.245 8.325 ;
        RECT 411.915 6.635 412.245 6.965 ;
        RECT 411.915 5.275 412.245 5.605 ;
        RECT 411.915 3.915 412.245 4.245 ;
        RECT 411.915 2.555 412.245 2.885 ;
        RECT 411.915 1.195 412.245 1.525 ;
        RECT 411.915 -0.165 412.245 0.165 ;
        RECT 411.92 -8.32 412.24 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 413.275 10.715 413.605 11.045 ;
        RECT 413.275 9.355 413.605 9.685 ;
        RECT 413.275 7.995 413.605 8.325 ;
        RECT 413.275 6.635 413.605 6.965 ;
        RECT 413.275 5.275 413.605 5.605 ;
        RECT 413.275 3.915 413.605 4.245 ;
        RECT 413.275 2.555 413.605 2.885 ;
        RECT 413.275 1.195 413.605 1.525 ;
        RECT 413.275 -0.165 413.605 0.165 ;
        RECT 413.28 -8.32 413.6 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 414.635 10.715 414.965 11.045 ;
        RECT 414.635 9.355 414.965 9.685 ;
        RECT 414.635 7.995 414.965 8.325 ;
        RECT 414.635 6.635 414.965 6.965 ;
        RECT 414.635 5.275 414.965 5.605 ;
        RECT 414.635 3.915 414.965 4.245 ;
        RECT 414.635 2.555 414.965 2.885 ;
        RECT 414.635 1.195 414.965 1.525 ;
        RECT 414.635 -0.165 414.965 0.165 ;
        RECT 414.64 -8.32 414.96 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 415.995 10.715 416.325 11.045 ;
        RECT 415.995 9.355 416.325 9.685 ;
        RECT 415.995 7.995 416.325 8.325 ;
        RECT 415.995 6.635 416.325 6.965 ;
        RECT 415.995 5.275 416.325 5.605 ;
        RECT 415.995 3.915 416.325 4.245 ;
        RECT 415.995 2.555 416.325 2.885 ;
        RECT 415.995 1.195 416.325 1.525 ;
        RECT 415.995 -0.165 416.325 0.165 ;
        RECT 416 -8.32 416.32 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 417.355 10.715 417.685 11.045 ;
        RECT 417.355 9.355 417.685 9.685 ;
        RECT 417.355 7.995 417.685 8.325 ;
        RECT 417.355 6.635 417.685 6.965 ;
        RECT 417.355 5.275 417.685 5.605 ;
        RECT 417.355 3.915 417.685 4.245 ;
        RECT 417.355 2.555 417.685 2.885 ;
        RECT 417.355 1.195 417.685 1.525 ;
        RECT 417.355 -0.165 417.685 0.165 ;
        RECT 417.36 -8.32 417.68 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 418.715 10.715 419.045 11.045 ;
        RECT 418.715 9.355 419.045 9.685 ;
        RECT 418.715 7.995 419.045 8.325 ;
        RECT 418.715 6.635 419.045 6.965 ;
        RECT 418.715 5.275 419.045 5.605 ;
        RECT 418.715 3.915 419.045 4.245 ;
        RECT 418.715 2.555 419.045 2.885 ;
        RECT 418.715 1.195 419.045 1.525 ;
        RECT 418.715 -0.165 419.045 0.165 ;
        RECT 418.72 -8.32 419.04 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 420.075 10.715 420.405 11.045 ;
        RECT 420.075 9.355 420.405 9.685 ;
        RECT 420.075 7.995 420.405 8.325 ;
        RECT 420.075 6.635 420.405 6.965 ;
        RECT 420.075 5.275 420.405 5.605 ;
        RECT 420.075 3.915 420.405 4.245 ;
        RECT 420.075 2.555 420.405 2.885 ;
        RECT 420.075 1.195 420.405 1.525 ;
        RECT 420.075 -0.165 420.405 0.165 ;
        RECT 420.08 -8.32 420.4 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 421.435 10.715 421.765 11.045 ;
        RECT 421.435 9.355 421.765 9.685 ;
        RECT 421.435 7.995 421.765 8.325 ;
        RECT 421.435 6.635 421.765 6.965 ;
        RECT 421.435 5.275 421.765 5.605 ;
        RECT 421.435 3.915 421.765 4.245 ;
        RECT 421.435 2.555 421.765 2.885 ;
        RECT 421.435 1.195 421.765 1.525 ;
        RECT 421.435 -0.165 421.765 0.165 ;
        RECT 421.44 -8.32 421.76 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 422.795 10.715 423.125 11.045 ;
        RECT 422.795 9.355 423.125 9.685 ;
        RECT 422.795 7.995 423.125 8.325 ;
        RECT 422.795 6.635 423.125 6.965 ;
        RECT 422.795 5.275 423.125 5.605 ;
        RECT 422.795 3.915 423.125 4.245 ;
        RECT 422.795 2.555 423.125 2.885 ;
        RECT 422.795 1.195 423.125 1.525 ;
        RECT 422.795 -0.165 423.125 0.165 ;
        RECT 422.8 -8.32 423.12 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 424.155 10.715 424.485 11.045 ;
        RECT 424.155 9.355 424.485 9.685 ;
        RECT 424.155 7.995 424.485 8.325 ;
        RECT 424.155 6.635 424.485 6.965 ;
        RECT 424.155 5.275 424.485 5.605 ;
        RECT 424.155 3.915 424.485 4.245 ;
        RECT 424.155 2.555 424.485 2.885 ;
        RECT 424.155 1.195 424.485 1.525 ;
        RECT 424.155 -0.165 424.485 0.165 ;
        RECT 424.16 -8.32 424.48 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 425.515 10.715 425.845 11.045 ;
        RECT 425.515 9.355 425.845 9.685 ;
        RECT 425.515 7.995 425.845 8.325 ;
        RECT 425.515 6.635 425.845 6.965 ;
        RECT 425.515 5.275 425.845 5.605 ;
        RECT 425.515 3.915 425.845 4.245 ;
        RECT 425.515 2.555 425.845 2.885 ;
        RECT 425.515 1.195 425.845 1.525 ;
        RECT 425.515 -0.165 425.845 0.165 ;
        RECT 425.52 -8.32 425.84 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 426.875 10.715 427.205 11.045 ;
        RECT 426.875 9.355 427.205 9.685 ;
        RECT 426.875 7.995 427.205 8.325 ;
        RECT 426.875 6.635 427.205 6.965 ;
        RECT 426.875 5.275 427.205 5.605 ;
        RECT 426.875 3.915 427.205 4.245 ;
        RECT 426.875 2.555 427.205 2.885 ;
        RECT 426.875 1.195 427.205 1.525 ;
        RECT 426.875 -0.165 427.205 0.165 ;
        RECT 426.88 -8.32 427.2 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 428.235 10.715 428.565 11.045 ;
        RECT 428.235 9.355 428.565 9.685 ;
        RECT 428.235 7.995 428.565 8.325 ;
        RECT 428.235 6.635 428.565 6.965 ;
        RECT 428.235 5.275 428.565 5.605 ;
        RECT 428.235 3.915 428.565 4.245 ;
        RECT 428.235 2.555 428.565 2.885 ;
        RECT 428.235 1.195 428.565 1.525 ;
        RECT 428.235 -0.165 428.565 0.165 ;
        RECT 428.24 -8.32 428.56 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 429.595 10.715 429.925 11.045 ;
        RECT 429.595 9.355 429.925 9.685 ;
        RECT 429.595 7.995 429.925 8.325 ;
        RECT 429.595 6.635 429.925 6.965 ;
        RECT 429.595 5.275 429.925 5.605 ;
        RECT 429.595 3.915 429.925 4.245 ;
        RECT 429.595 2.555 429.925 2.885 ;
        RECT 429.595 1.195 429.925 1.525 ;
        RECT 429.595 -0.165 429.925 0.165 ;
        RECT 429.6 -8.32 429.92 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 430.955 10.715 431.285 11.045 ;
        RECT 430.955 9.355 431.285 9.685 ;
        RECT 430.955 7.995 431.285 8.325 ;
        RECT 430.955 6.635 431.285 6.965 ;
        RECT 430.955 5.275 431.285 5.605 ;
        RECT 430.955 3.915 431.285 4.245 ;
        RECT 430.955 2.555 431.285 2.885 ;
        RECT 430.955 1.195 431.285 1.525 ;
        RECT 430.955 -0.165 431.285 0.165 ;
        RECT 430.96 -8.32 431.28 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 432.315 10.715 432.645 11.045 ;
        RECT 432.315 9.355 432.645 9.685 ;
        RECT 432.315 7.995 432.645 8.325 ;
        RECT 432.315 6.635 432.645 6.965 ;
        RECT 432.315 5.275 432.645 5.605 ;
        RECT 432.315 3.915 432.645 4.245 ;
        RECT 432.315 2.555 432.645 2.885 ;
        RECT 432.315 1.195 432.645 1.525 ;
        RECT 432.315 -0.165 432.645 0.165 ;
        RECT 432.32 -8.32 432.64 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 433.675 10.715 434.005 11.045 ;
        RECT 433.675 9.355 434.005 9.685 ;
        RECT 433.675 7.995 434.005 8.325 ;
        RECT 433.675 6.635 434.005 6.965 ;
        RECT 433.675 5.275 434.005 5.605 ;
        RECT 433.675 3.915 434.005 4.245 ;
        RECT 433.675 2.555 434.005 2.885 ;
        RECT 433.675 1.195 434.005 1.525 ;
        RECT 433.675 -0.165 434.005 0.165 ;
        RECT 433.68 -8.32 434 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 435.035 10.715 435.365 11.045 ;
        RECT 435.035 9.355 435.365 9.685 ;
        RECT 435.035 7.995 435.365 8.325 ;
        RECT 435.035 6.635 435.365 6.965 ;
        RECT 435.035 5.275 435.365 5.605 ;
        RECT 435.035 3.915 435.365 4.245 ;
        RECT 435.035 2.555 435.365 2.885 ;
        RECT 435.035 1.195 435.365 1.525 ;
        RECT 435.035 -0.165 435.365 0.165 ;
        RECT 435.04 -8.32 435.36 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 436.395 10.715 436.725 11.045 ;
        RECT 436.395 9.355 436.725 9.685 ;
        RECT 436.395 7.995 436.725 8.325 ;
        RECT 436.395 6.635 436.725 6.965 ;
        RECT 436.395 5.275 436.725 5.605 ;
        RECT 436.395 3.915 436.725 4.245 ;
        RECT 436.395 2.555 436.725 2.885 ;
        RECT 436.395 1.195 436.725 1.525 ;
        RECT 436.395 -0.165 436.725 0.165 ;
        RECT 436.4 -8.32 436.72 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 437.755 10.715 438.085 11.045 ;
        RECT 437.755 9.355 438.085 9.685 ;
        RECT 437.755 7.995 438.085 8.325 ;
        RECT 437.755 6.635 438.085 6.965 ;
        RECT 437.755 5.275 438.085 5.605 ;
        RECT 437.755 3.915 438.085 4.245 ;
        RECT 437.755 2.555 438.085 2.885 ;
        RECT 437.755 1.195 438.085 1.525 ;
        RECT 437.755 -0.165 438.085 0.165 ;
        RECT 437.76 -8.32 438.08 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 439.115 10.715 439.445 11.045 ;
        RECT 439.115 9.355 439.445 9.685 ;
        RECT 439.115 7.995 439.445 8.325 ;
        RECT 439.115 6.635 439.445 6.965 ;
        RECT 439.115 5.275 439.445 5.605 ;
        RECT 439.115 3.915 439.445 4.245 ;
        RECT 439.115 2.555 439.445 2.885 ;
        RECT 439.115 1.195 439.445 1.525 ;
        RECT 439.115 -0.165 439.445 0.165 ;
        RECT 439.12 -8.32 439.44 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 440.475 10.715 440.805 11.045 ;
        RECT 440.475 9.355 440.805 9.685 ;
        RECT 440.475 7.995 440.805 8.325 ;
        RECT 440.475 6.635 440.805 6.965 ;
        RECT 440.475 5.275 440.805 5.605 ;
        RECT 440.475 3.915 440.805 4.245 ;
        RECT 440.475 2.555 440.805 2.885 ;
        RECT 440.475 1.195 440.805 1.525 ;
        RECT 440.475 -0.165 440.805 0.165 ;
        RECT 440.48 -8.32 440.8 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 441.835 10.715 442.165 11.045 ;
        RECT 441.835 9.355 442.165 9.685 ;
        RECT 441.835 7.995 442.165 8.325 ;
        RECT 441.835 6.635 442.165 6.965 ;
        RECT 441.835 5.275 442.165 5.605 ;
        RECT 441.835 3.915 442.165 4.245 ;
        RECT 441.835 2.555 442.165 2.885 ;
        RECT 441.835 1.195 442.165 1.525 ;
        RECT 441.835 -0.165 442.165 0.165 ;
        RECT 441.84 -8.32 442.16 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 443.195 10.715 443.525 11.045 ;
        RECT 443.195 9.355 443.525 9.685 ;
        RECT 443.195 7.995 443.525 8.325 ;
        RECT 443.195 6.635 443.525 6.965 ;
        RECT 443.195 5.275 443.525 5.605 ;
        RECT 443.195 3.915 443.525 4.245 ;
        RECT 443.195 2.555 443.525 2.885 ;
        RECT 443.195 1.195 443.525 1.525 ;
        RECT 443.195 -0.165 443.525 0.165 ;
        RECT 443.2 -8.32 443.52 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 444.555 10.715 444.885 11.045 ;
        RECT 444.555 9.355 444.885 9.685 ;
        RECT 444.555 7.995 444.885 8.325 ;
        RECT 444.555 6.635 444.885 6.965 ;
        RECT 444.555 5.275 444.885 5.605 ;
        RECT 444.555 3.915 444.885 4.245 ;
        RECT 444.555 2.555 444.885 2.885 ;
        RECT 444.555 1.195 444.885 1.525 ;
        RECT 444.555 -0.165 444.885 0.165 ;
        RECT 444.56 -8.32 444.88 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 445.915 10.715 446.245 11.045 ;
        RECT 445.915 9.355 446.245 9.685 ;
        RECT 445.915 7.995 446.245 8.325 ;
        RECT 445.915 6.635 446.245 6.965 ;
        RECT 445.915 5.275 446.245 5.605 ;
        RECT 445.915 3.915 446.245 4.245 ;
        RECT 445.915 2.555 446.245 2.885 ;
        RECT 445.915 1.195 446.245 1.525 ;
        RECT 445.915 -0.165 446.245 0.165 ;
        RECT 445.92 -8.32 446.24 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 447.275 10.715 447.605 11.045 ;
        RECT 447.275 9.355 447.605 9.685 ;
        RECT 447.275 7.995 447.605 8.325 ;
        RECT 447.275 6.635 447.605 6.965 ;
        RECT 447.275 5.275 447.605 5.605 ;
        RECT 447.275 3.915 447.605 4.245 ;
        RECT 447.275 2.555 447.605 2.885 ;
        RECT 447.275 1.195 447.605 1.525 ;
        RECT 447.275 -0.165 447.605 0.165 ;
        RECT 447.28 -8.32 447.6 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 448.635 10.715 448.965 11.045 ;
        RECT 448.635 9.355 448.965 9.685 ;
        RECT 448.635 7.995 448.965 8.325 ;
        RECT 448.635 6.635 448.965 6.965 ;
        RECT 448.635 5.275 448.965 5.605 ;
        RECT 448.635 3.915 448.965 4.245 ;
        RECT 448.635 2.555 448.965 2.885 ;
        RECT 448.635 1.195 448.965 1.525 ;
        RECT 448.635 -0.165 448.965 0.165 ;
        RECT 448.64 -8.32 448.96 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 449.995 10.715 450.325 11.045 ;
        RECT 449.995 9.355 450.325 9.685 ;
        RECT 449.995 7.995 450.325 8.325 ;
        RECT 449.995 6.635 450.325 6.965 ;
        RECT 449.995 5.275 450.325 5.605 ;
        RECT 449.995 3.915 450.325 4.245 ;
        RECT 449.995 2.555 450.325 2.885 ;
        RECT 449.995 1.195 450.325 1.525 ;
        RECT 449.995 -0.165 450.325 0.165 ;
        RECT 450 -8.32 450.32 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 451.355 10.715 451.685 11.045 ;
        RECT 451.355 9.355 451.685 9.685 ;
        RECT 451.355 7.995 451.685 8.325 ;
        RECT 451.355 6.635 451.685 6.965 ;
        RECT 451.355 5.275 451.685 5.605 ;
        RECT 451.355 3.915 451.685 4.245 ;
        RECT 451.355 2.555 451.685 2.885 ;
        RECT 451.355 1.195 451.685 1.525 ;
        RECT 451.355 -0.165 451.685 0.165 ;
        RECT 451.36 -8.32 451.68 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 452.715 10.715 453.045 11.045 ;
        RECT 452.715 9.355 453.045 9.685 ;
        RECT 452.715 7.995 453.045 8.325 ;
        RECT 452.715 6.635 453.045 6.965 ;
        RECT 452.715 5.275 453.045 5.605 ;
        RECT 452.715 3.915 453.045 4.245 ;
        RECT 452.715 2.555 453.045 2.885 ;
        RECT 452.715 1.195 453.045 1.525 ;
        RECT 452.715 -0.165 453.045 0.165 ;
        RECT 452.72 -8.32 453.04 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 454.075 10.715 454.405 11.045 ;
        RECT 454.075 9.355 454.405 9.685 ;
        RECT 454.075 7.995 454.405 8.325 ;
        RECT 454.075 6.635 454.405 6.965 ;
        RECT 454.075 5.275 454.405 5.605 ;
        RECT 454.075 3.915 454.405 4.245 ;
        RECT 454.075 2.555 454.405 2.885 ;
        RECT 454.075 1.195 454.405 1.525 ;
        RECT 454.075 -0.165 454.405 0.165 ;
        RECT 454.08 -8.32 454.4 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 455.435 10.715 455.765 11.045 ;
        RECT 455.435 9.355 455.765 9.685 ;
        RECT 455.435 7.995 455.765 8.325 ;
        RECT 455.435 6.635 455.765 6.965 ;
        RECT 455.435 5.275 455.765 5.605 ;
        RECT 455.435 3.915 455.765 4.245 ;
        RECT 455.435 2.555 455.765 2.885 ;
        RECT 455.435 1.195 455.765 1.525 ;
        RECT 455.435 -0.165 455.765 0.165 ;
        RECT 455.44 -8.32 455.76 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 456.795 10.715 457.125 11.045 ;
        RECT 456.795 9.355 457.125 9.685 ;
        RECT 456.795 7.995 457.125 8.325 ;
        RECT 456.795 6.635 457.125 6.965 ;
        RECT 456.795 5.275 457.125 5.605 ;
        RECT 456.795 3.915 457.125 4.245 ;
        RECT 456.795 2.555 457.125 2.885 ;
        RECT 456.795 1.195 457.125 1.525 ;
        RECT 456.795 -0.165 457.125 0.165 ;
        RECT 456.8 -8.32 457.12 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 458.155 10.715 458.485 11.045 ;
        RECT 458.155 9.355 458.485 9.685 ;
        RECT 458.155 7.995 458.485 8.325 ;
        RECT 458.155 6.635 458.485 6.965 ;
        RECT 458.155 5.275 458.485 5.605 ;
        RECT 458.155 3.915 458.485 4.245 ;
        RECT 458.155 2.555 458.485 2.885 ;
        RECT 458.155 1.195 458.485 1.525 ;
        RECT 458.155 -0.165 458.485 0.165 ;
        RECT 458.16 -8.32 458.48 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 459.515 10.715 459.845 11.045 ;
        RECT 459.515 9.355 459.845 9.685 ;
        RECT 459.515 7.995 459.845 8.325 ;
        RECT 459.515 6.635 459.845 6.965 ;
        RECT 459.515 5.275 459.845 5.605 ;
        RECT 459.515 3.915 459.845 4.245 ;
        RECT 459.515 2.555 459.845 2.885 ;
        RECT 459.515 1.195 459.845 1.525 ;
        RECT 459.515 -0.165 459.845 0.165 ;
        RECT 459.52 -8.32 459.84 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 460.875 10.715 461.205 11.045 ;
        RECT 460.875 9.355 461.205 9.685 ;
        RECT 460.875 7.995 461.205 8.325 ;
        RECT 460.875 6.635 461.205 6.965 ;
        RECT 460.875 5.275 461.205 5.605 ;
        RECT 460.875 3.915 461.205 4.245 ;
        RECT 460.875 2.555 461.205 2.885 ;
        RECT 460.875 1.195 461.205 1.525 ;
        RECT 460.875 -0.165 461.205 0.165 ;
        RECT 460.88 -8.32 461.2 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 462.235 10.715 462.565 11.045 ;
        RECT 462.235 9.355 462.565 9.685 ;
        RECT 462.235 7.995 462.565 8.325 ;
        RECT 462.235 6.635 462.565 6.965 ;
        RECT 462.235 5.275 462.565 5.605 ;
        RECT 462.235 3.915 462.565 4.245 ;
        RECT 462.235 2.555 462.565 2.885 ;
        RECT 462.235 1.195 462.565 1.525 ;
        RECT 462.235 -0.165 462.565 0.165 ;
        RECT 462.24 -8.32 462.56 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 463.595 10.715 463.925 11.045 ;
        RECT 463.595 9.355 463.925 9.685 ;
        RECT 463.595 7.995 463.925 8.325 ;
        RECT 463.595 6.635 463.925 6.965 ;
        RECT 463.595 5.275 463.925 5.605 ;
        RECT 463.595 3.915 463.925 4.245 ;
        RECT 463.595 2.555 463.925 2.885 ;
        RECT 463.595 1.195 463.925 1.525 ;
        RECT 463.595 -0.165 463.925 0.165 ;
        RECT 463.6 -8.32 463.92 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 464.955 10.715 465.285 11.045 ;
        RECT 464.955 9.355 465.285 9.685 ;
        RECT 464.955 7.995 465.285 8.325 ;
        RECT 464.955 6.635 465.285 6.965 ;
        RECT 464.955 5.275 465.285 5.605 ;
        RECT 464.955 3.915 465.285 4.245 ;
        RECT 464.955 2.555 465.285 2.885 ;
        RECT 464.955 1.195 465.285 1.525 ;
        RECT 464.955 -0.165 465.285 0.165 ;
        RECT 464.96 -8.32 465.28 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 466.315 10.715 466.645 11.045 ;
        RECT 466.315 9.355 466.645 9.685 ;
        RECT 466.315 7.995 466.645 8.325 ;
        RECT 466.315 6.635 466.645 6.965 ;
        RECT 466.315 5.275 466.645 5.605 ;
        RECT 466.315 3.915 466.645 4.245 ;
        RECT 466.315 2.555 466.645 2.885 ;
        RECT 466.315 1.195 466.645 1.525 ;
        RECT 466.315 -0.165 466.645 0.165 ;
        RECT 466.32 -8.32 466.64 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 467.675 10.715 468.005 11.045 ;
        RECT 467.675 9.355 468.005 9.685 ;
        RECT 467.675 7.995 468.005 8.325 ;
        RECT 467.675 6.635 468.005 6.965 ;
        RECT 467.675 5.275 468.005 5.605 ;
        RECT 467.675 3.915 468.005 4.245 ;
        RECT 467.675 2.555 468.005 2.885 ;
        RECT 467.675 1.195 468.005 1.525 ;
        RECT 467.675 -0.165 468.005 0.165 ;
        RECT 467.68 -8.32 468 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 469.035 10.715 469.365 11.045 ;
        RECT 469.035 9.355 469.365 9.685 ;
        RECT 469.035 7.995 469.365 8.325 ;
        RECT 469.035 6.635 469.365 6.965 ;
        RECT 469.035 5.275 469.365 5.605 ;
        RECT 469.035 3.915 469.365 4.245 ;
        RECT 469.035 2.555 469.365 2.885 ;
        RECT 469.035 1.195 469.365 1.525 ;
        RECT 469.035 -0.165 469.365 0.165 ;
        RECT 469.04 -8.32 469.36 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 470.395 10.715 470.725 11.045 ;
        RECT 470.395 9.355 470.725 9.685 ;
        RECT 470.395 7.995 470.725 8.325 ;
        RECT 470.395 6.635 470.725 6.965 ;
        RECT 470.395 5.275 470.725 5.605 ;
        RECT 470.395 3.915 470.725 4.245 ;
        RECT 470.395 2.555 470.725 2.885 ;
        RECT 470.395 1.195 470.725 1.525 ;
        RECT 470.395 -0.165 470.725 0.165 ;
        RECT 470.4 -8.32 470.72 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 471.755 10.715 472.085 11.045 ;
        RECT 471.755 9.355 472.085 9.685 ;
        RECT 471.755 7.995 472.085 8.325 ;
        RECT 471.755 6.635 472.085 6.965 ;
        RECT 471.755 5.275 472.085 5.605 ;
        RECT 471.755 3.915 472.085 4.245 ;
        RECT 471.755 2.555 472.085 2.885 ;
        RECT 471.755 1.195 472.085 1.525 ;
        RECT 471.755 -0.165 472.085 0.165 ;
        RECT 471.76 -8.32 472.08 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 473.115 10.715 473.445 11.045 ;
        RECT 473.115 9.355 473.445 9.685 ;
        RECT 473.115 7.995 473.445 8.325 ;
        RECT 473.115 6.635 473.445 6.965 ;
        RECT 473.115 5.275 473.445 5.605 ;
        RECT 473.115 3.915 473.445 4.245 ;
        RECT 473.115 2.555 473.445 2.885 ;
        RECT 473.115 1.195 473.445 1.525 ;
        RECT 473.115 -0.165 473.445 0.165 ;
        RECT 473.12 -8.32 473.44 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 474.475 10.715 474.805 11.045 ;
        RECT 474.475 9.355 474.805 9.685 ;
        RECT 474.475 7.995 474.805 8.325 ;
        RECT 474.475 6.635 474.805 6.965 ;
        RECT 474.475 5.275 474.805 5.605 ;
        RECT 474.475 3.915 474.805 4.245 ;
        RECT 474.475 2.555 474.805 2.885 ;
        RECT 474.475 1.195 474.805 1.525 ;
        RECT 474.475 -0.165 474.805 0.165 ;
        RECT 474.48 -8.32 474.8 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 475.835 10.715 476.165 11.045 ;
        RECT 475.835 9.355 476.165 9.685 ;
        RECT 475.835 7.995 476.165 8.325 ;
        RECT 475.835 6.635 476.165 6.965 ;
        RECT 475.835 5.275 476.165 5.605 ;
        RECT 475.835 3.915 476.165 4.245 ;
        RECT 475.835 2.555 476.165 2.885 ;
        RECT 475.835 1.195 476.165 1.525 ;
        RECT 475.835 -0.165 476.165 0.165 ;
        RECT 475.84 -8.32 476.16 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 477.195 10.715 477.525 11.045 ;
        RECT 477.195 9.355 477.525 9.685 ;
        RECT 477.195 7.995 477.525 8.325 ;
        RECT 477.195 6.635 477.525 6.965 ;
        RECT 477.195 5.275 477.525 5.605 ;
        RECT 477.195 3.915 477.525 4.245 ;
        RECT 477.195 2.555 477.525 2.885 ;
        RECT 477.195 1.195 477.525 1.525 ;
        RECT 477.195 -0.165 477.525 0.165 ;
        RECT 477.2 -8.32 477.52 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 478.555 10.715 478.885 11.045 ;
        RECT 478.555 9.355 478.885 9.685 ;
        RECT 478.555 7.995 478.885 8.325 ;
        RECT 478.555 6.635 478.885 6.965 ;
        RECT 478.555 5.275 478.885 5.605 ;
        RECT 478.555 3.915 478.885 4.245 ;
        RECT 478.555 2.555 478.885 2.885 ;
        RECT 478.555 1.195 478.885 1.525 ;
        RECT 478.555 -0.165 478.885 0.165 ;
        RECT 478.56 -8.32 478.88 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 479.915 10.715 480.245 11.045 ;
        RECT 479.915 9.355 480.245 9.685 ;
        RECT 479.915 7.995 480.245 8.325 ;
        RECT 479.915 6.635 480.245 6.965 ;
        RECT 479.915 5.275 480.245 5.605 ;
        RECT 479.915 3.915 480.245 4.245 ;
        RECT 479.915 2.555 480.245 2.885 ;
        RECT 479.915 1.195 480.245 1.525 ;
        RECT 479.915 -0.165 480.245 0.165 ;
        RECT 479.92 -8.32 480.24 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 481.275 10.715 481.605 11.045 ;
        RECT 481.275 9.355 481.605 9.685 ;
        RECT 481.275 7.995 481.605 8.325 ;
        RECT 481.275 6.635 481.605 6.965 ;
        RECT 481.275 5.275 481.605 5.605 ;
        RECT 481.275 3.915 481.605 4.245 ;
        RECT 481.275 2.555 481.605 2.885 ;
        RECT 481.275 1.195 481.605 1.525 ;
        RECT 481.275 -0.165 481.605 0.165 ;
        RECT 481.28 -8.32 481.6 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 482.635 10.715 482.965 11.045 ;
        RECT 482.635 9.355 482.965 9.685 ;
        RECT 482.635 7.995 482.965 8.325 ;
        RECT 482.635 6.635 482.965 6.965 ;
        RECT 482.635 5.275 482.965 5.605 ;
        RECT 482.635 3.915 482.965 4.245 ;
        RECT 482.635 2.555 482.965 2.885 ;
        RECT 482.635 1.195 482.965 1.525 ;
        RECT 482.635 -0.165 482.965 0.165 ;
        RECT 482.64 -8.32 482.96 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 483.995 10.715 484.325 11.045 ;
        RECT 483.995 9.355 484.325 9.685 ;
        RECT 483.995 7.995 484.325 8.325 ;
        RECT 483.995 6.635 484.325 6.965 ;
        RECT 483.995 5.275 484.325 5.605 ;
        RECT 483.995 3.915 484.325 4.245 ;
        RECT 483.995 2.555 484.325 2.885 ;
        RECT 483.995 1.195 484.325 1.525 ;
        RECT 483.995 -0.165 484.325 0.165 ;
        RECT 484 -8.32 484.32 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 485.355 10.715 485.685 11.045 ;
        RECT 485.355 9.355 485.685 9.685 ;
        RECT 485.355 7.995 485.685 8.325 ;
        RECT 485.355 6.635 485.685 6.965 ;
        RECT 485.355 5.275 485.685 5.605 ;
        RECT 485.355 3.915 485.685 4.245 ;
        RECT 485.355 2.555 485.685 2.885 ;
        RECT 485.355 1.195 485.685 1.525 ;
        RECT 485.355 -0.165 485.685 0.165 ;
        RECT 485.36 -8.32 485.68 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 486.715 10.715 487.045 11.045 ;
        RECT 486.715 9.355 487.045 9.685 ;
        RECT 486.715 7.995 487.045 8.325 ;
        RECT 486.715 6.635 487.045 6.965 ;
        RECT 486.715 5.275 487.045 5.605 ;
        RECT 486.715 3.915 487.045 4.245 ;
        RECT 486.715 2.555 487.045 2.885 ;
        RECT 486.715 1.195 487.045 1.525 ;
        RECT 486.715 -0.165 487.045 0.165 ;
        RECT 486.72 -8.32 487.04 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 488.075 10.715 488.405 11.045 ;
        RECT 488.075 9.355 488.405 9.685 ;
        RECT 488.075 7.995 488.405 8.325 ;
        RECT 488.075 6.635 488.405 6.965 ;
        RECT 488.075 5.275 488.405 5.605 ;
        RECT 488.075 3.915 488.405 4.245 ;
        RECT 488.075 2.555 488.405 2.885 ;
        RECT 488.075 1.195 488.405 1.525 ;
        RECT 488.075 -0.165 488.405 0.165 ;
        RECT 488.08 -8.32 488.4 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 489.435 10.715 489.765 11.045 ;
        RECT 489.435 9.355 489.765 9.685 ;
        RECT 489.435 7.995 489.765 8.325 ;
        RECT 489.435 6.635 489.765 6.965 ;
        RECT 489.435 5.275 489.765 5.605 ;
        RECT 489.435 3.915 489.765 4.245 ;
        RECT 489.435 2.555 489.765 2.885 ;
        RECT 489.435 1.195 489.765 1.525 ;
        RECT 489.435 -0.165 489.765 0.165 ;
        RECT 489.44 -8.32 489.76 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 490.795 10.715 491.125 11.045 ;
        RECT 490.795 9.355 491.125 9.685 ;
        RECT 490.795 7.995 491.125 8.325 ;
        RECT 490.795 6.635 491.125 6.965 ;
        RECT 490.795 5.275 491.125 5.605 ;
        RECT 490.795 3.915 491.125 4.245 ;
        RECT 490.795 2.555 491.125 2.885 ;
        RECT 490.795 1.195 491.125 1.525 ;
        RECT 490.795 -0.165 491.125 0.165 ;
        RECT 490.8 -8.32 491.12 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 492.155 10.715 492.485 11.045 ;
        RECT 492.155 9.355 492.485 9.685 ;
        RECT 492.155 7.995 492.485 8.325 ;
        RECT 492.155 6.635 492.485 6.965 ;
        RECT 492.155 5.275 492.485 5.605 ;
        RECT 492.155 3.915 492.485 4.245 ;
        RECT 492.155 2.555 492.485 2.885 ;
        RECT 492.155 1.195 492.485 1.525 ;
        RECT 492.155 -0.165 492.485 0.165 ;
        RECT 492.16 -8.32 492.48 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 493.515 10.715 493.845 11.045 ;
        RECT 493.515 9.355 493.845 9.685 ;
        RECT 493.515 7.995 493.845 8.325 ;
        RECT 493.515 6.635 493.845 6.965 ;
        RECT 493.515 5.275 493.845 5.605 ;
        RECT 493.515 3.915 493.845 4.245 ;
        RECT 493.515 2.555 493.845 2.885 ;
        RECT 493.515 1.195 493.845 1.525 ;
        RECT 493.515 -0.165 493.845 0.165 ;
        RECT 493.52 -8.32 493.84 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 494.875 10.715 495.205 11.045 ;
        RECT 494.875 9.355 495.205 9.685 ;
        RECT 494.875 7.995 495.205 8.325 ;
        RECT 494.875 6.635 495.205 6.965 ;
        RECT 494.875 5.275 495.205 5.605 ;
        RECT 494.875 3.915 495.205 4.245 ;
        RECT 494.875 2.555 495.205 2.885 ;
        RECT 494.875 1.195 495.205 1.525 ;
        RECT 494.875 -0.165 495.205 0.165 ;
        RECT 494.88 -8.32 495.2 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 496.235 10.715 496.565 11.045 ;
        RECT 496.235 9.355 496.565 9.685 ;
        RECT 496.235 7.995 496.565 8.325 ;
        RECT 496.235 6.635 496.565 6.965 ;
        RECT 496.235 5.275 496.565 5.605 ;
        RECT 496.235 3.915 496.565 4.245 ;
        RECT 496.235 2.555 496.565 2.885 ;
        RECT 496.235 1.195 496.565 1.525 ;
        RECT 496.235 -0.165 496.565 0.165 ;
        RECT 496.24 -8.32 496.56 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 497.595 9.355 497.925 9.685 ;
        RECT 497.595 7.995 497.925 8.325 ;
        RECT 497.595 6.635 497.925 6.965 ;
        RECT 497.595 5.275 497.925 5.605 ;
        RECT 497.595 3.915 497.925 4.245 ;
        RECT 497.595 2.555 497.925 2.885 ;
        RECT 497.595 1.195 497.925 1.525 ;
        RECT 497.595 -0.165 497.925 0.165 ;
        RECT 497.6 -8.32 497.92 15.8 ;
        RECT 497.595 10.715 497.925 11.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.955 10.715 227.285 11.045 ;
        RECT 226.955 9.355 227.285 9.685 ;
        RECT 226.955 7.995 227.285 8.325 ;
        RECT 226.955 6.635 227.285 6.965 ;
        RECT 226.955 5.275 227.285 5.605 ;
        RECT 226.955 3.915 227.285 4.245 ;
        RECT 226.955 2.555 227.285 2.885 ;
        RECT 226.955 1.195 227.285 1.525 ;
        RECT 226.955 -0.165 227.285 0.165 ;
        RECT 226.96 -8.32 227.28 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.315 10.715 228.645 11.045 ;
        RECT 228.315 9.355 228.645 9.685 ;
        RECT 228.315 7.995 228.645 8.325 ;
        RECT 228.315 6.635 228.645 6.965 ;
        RECT 228.315 5.275 228.645 5.605 ;
        RECT 228.315 3.915 228.645 4.245 ;
        RECT 228.315 2.555 228.645 2.885 ;
        RECT 228.315 1.195 228.645 1.525 ;
        RECT 228.315 -0.165 228.645 0.165 ;
        RECT 228.32 -8.32 228.64 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 229.675 10.715 230.005 11.045 ;
        RECT 229.675 9.355 230.005 9.685 ;
        RECT 229.675 7.995 230.005 8.325 ;
        RECT 229.675 6.635 230.005 6.965 ;
        RECT 229.675 5.275 230.005 5.605 ;
        RECT 229.675 3.915 230.005 4.245 ;
        RECT 229.675 2.555 230.005 2.885 ;
        RECT 229.675 1.195 230.005 1.525 ;
        RECT 229.675 -0.165 230.005 0.165 ;
        RECT 229.68 -8.32 230 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 231.035 10.715 231.365 11.045 ;
        RECT 231.035 9.355 231.365 9.685 ;
        RECT 231.035 7.995 231.365 8.325 ;
        RECT 231.035 6.635 231.365 6.965 ;
        RECT 231.035 5.275 231.365 5.605 ;
        RECT 231.035 3.915 231.365 4.245 ;
        RECT 231.035 2.555 231.365 2.885 ;
        RECT 231.035 1.195 231.365 1.525 ;
        RECT 231.035 -0.165 231.365 0.165 ;
        RECT 231.04 -8.32 231.36 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 232.395 10.715 232.725 11.045 ;
        RECT 232.395 9.355 232.725 9.685 ;
        RECT 232.395 7.995 232.725 8.325 ;
        RECT 232.395 6.635 232.725 6.965 ;
        RECT 232.395 5.275 232.725 5.605 ;
        RECT 232.395 3.915 232.725 4.245 ;
        RECT 232.395 2.555 232.725 2.885 ;
        RECT 232.395 1.195 232.725 1.525 ;
        RECT 232.395 -0.165 232.725 0.165 ;
        RECT 232.4 -8.32 232.72 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.755 10.715 234.085 11.045 ;
        RECT 233.755 9.355 234.085 9.685 ;
        RECT 233.755 7.995 234.085 8.325 ;
        RECT 233.755 6.635 234.085 6.965 ;
        RECT 233.755 5.275 234.085 5.605 ;
        RECT 233.755 3.915 234.085 4.245 ;
        RECT 233.755 2.555 234.085 2.885 ;
        RECT 233.755 1.195 234.085 1.525 ;
        RECT 233.755 -0.165 234.085 0.165 ;
        RECT 233.76 -8.32 234.08 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 235.115 10.715 235.445 11.045 ;
        RECT 235.115 9.355 235.445 9.685 ;
        RECT 235.115 7.995 235.445 8.325 ;
        RECT 235.115 6.635 235.445 6.965 ;
        RECT 235.115 5.275 235.445 5.605 ;
        RECT 235.115 3.915 235.445 4.245 ;
        RECT 235.115 2.555 235.445 2.885 ;
        RECT 235.115 1.195 235.445 1.525 ;
        RECT 235.115 -0.165 235.445 0.165 ;
        RECT 235.12 -8.32 235.44 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 236.475 10.715 236.805 11.045 ;
        RECT 236.475 9.355 236.805 9.685 ;
        RECT 236.475 7.995 236.805 8.325 ;
        RECT 236.475 6.635 236.805 6.965 ;
        RECT 236.475 5.275 236.805 5.605 ;
        RECT 236.475 3.915 236.805 4.245 ;
        RECT 236.475 2.555 236.805 2.885 ;
        RECT 236.475 1.195 236.805 1.525 ;
        RECT 236.475 -0.165 236.805 0.165 ;
        RECT 236.48 -8.32 236.8 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 237.835 10.715 238.165 11.045 ;
        RECT 237.835 9.355 238.165 9.685 ;
        RECT 237.835 7.995 238.165 8.325 ;
        RECT 237.835 6.635 238.165 6.965 ;
        RECT 237.835 5.275 238.165 5.605 ;
        RECT 237.835 3.915 238.165 4.245 ;
        RECT 237.835 2.555 238.165 2.885 ;
        RECT 237.835 1.195 238.165 1.525 ;
        RECT 237.835 -0.165 238.165 0.165 ;
        RECT 237.84 -8.32 238.16 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.195 10.715 239.525 11.045 ;
        RECT 239.195 9.355 239.525 9.685 ;
        RECT 239.195 7.995 239.525 8.325 ;
        RECT 239.195 6.635 239.525 6.965 ;
        RECT 239.195 5.275 239.525 5.605 ;
        RECT 239.195 3.915 239.525 4.245 ;
        RECT 239.195 2.555 239.525 2.885 ;
        RECT 239.195 1.195 239.525 1.525 ;
        RECT 239.195 -0.165 239.525 0.165 ;
        RECT 239.2 -8.32 239.52 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 240.555 10.715 240.885 11.045 ;
        RECT 240.555 9.355 240.885 9.685 ;
        RECT 240.555 7.995 240.885 8.325 ;
        RECT 240.555 6.635 240.885 6.965 ;
        RECT 240.555 5.275 240.885 5.605 ;
        RECT 240.555 3.915 240.885 4.245 ;
        RECT 240.555 2.555 240.885 2.885 ;
        RECT 240.555 1.195 240.885 1.525 ;
        RECT 240.555 -0.165 240.885 0.165 ;
        RECT 240.56 -8.32 240.88 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 241.915 10.715 242.245 11.045 ;
        RECT 241.915 9.355 242.245 9.685 ;
        RECT 241.915 7.995 242.245 8.325 ;
        RECT 241.915 6.635 242.245 6.965 ;
        RECT 241.915 5.275 242.245 5.605 ;
        RECT 241.915 3.915 242.245 4.245 ;
        RECT 241.915 2.555 242.245 2.885 ;
        RECT 241.915 1.195 242.245 1.525 ;
        RECT 241.915 -0.165 242.245 0.165 ;
        RECT 241.92 -8.32 242.24 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 243.275 10.715 243.605 11.045 ;
        RECT 243.275 9.355 243.605 9.685 ;
        RECT 243.275 7.995 243.605 8.325 ;
        RECT 243.275 6.635 243.605 6.965 ;
        RECT 243.275 5.275 243.605 5.605 ;
        RECT 243.275 3.915 243.605 4.245 ;
        RECT 243.275 2.555 243.605 2.885 ;
        RECT 243.275 1.195 243.605 1.525 ;
        RECT 243.275 -0.165 243.605 0.165 ;
        RECT 243.28 -8.32 243.6 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 244.635 10.715 244.965 11.045 ;
        RECT 244.635 9.355 244.965 9.685 ;
        RECT 244.635 7.995 244.965 8.325 ;
        RECT 244.635 6.635 244.965 6.965 ;
        RECT 244.635 5.275 244.965 5.605 ;
        RECT 244.635 3.915 244.965 4.245 ;
        RECT 244.635 2.555 244.965 2.885 ;
        RECT 244.635 1.195 244.965 1.525 ;
        RECT 244.635 -0.165 244.965 0.165 ;
        RECT 244.64 -8.32 244.96 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 245.995 10.715 246.325 11.045 ;
        RECT 245.995 9.355 246.325 9.685 ;
        RECT 245.995 7.995 246.325 8.325 ;
        RECT 245.995 6.635 246.325 6.965 ;
        RECT 245.995 5.275 246.325 5.605 ;
        RECT 245.995 3.915 246.325 4.245 ;
        RECT 245.995 2.555 246.325 2.885 ;
        RECT 245.995 1.195 246.325 1.525 ;
        RECT 245.995 -0.165 246.325 0.165 ;
        RECT 246 -8.32 246.32 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 247.355 10.715 247.685 11.045 ;
        RECT 247.355 9.355 247.685 9.685 ;
        RECT 247.355 7.995 247.685 8.325 ;
        RECT 247.355 6.635 247.685 6.965 ;
        RECT 247.355 5.275 247.685 5.605 ;
        RECT 247.355 3.915 247.685 4.245 ;
        RECT 247.355 2.555 247.685 2.885 ;
        RECT 247.355 1.195 247.685 1.525 ;
        RECT 247.355 -0.165 247.685 0.165 ;
        RECT 247.36 -8.32 247.68 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.715 10.715 249.045 11.045 ;
        RECT 248.715 9.355 249.045 9.685 ;
        RECT 248.715 7.995 249.045 8.325 ;
        RECT 248.715 6.635 249.045 6.965 ;
        RECT 248.715 5.275 249.045 5.605 ;
        RECT 248.715 3.915 249.045 4.245 ;
        RECT 248.715 2.555 249.045 2.885 ;
        RECT 248.715 1.195 249.045 1.525 ;
        RECT 248.715 -0.165 249.045 0.165 ;
        RECT 248.72 -8.32 249.04 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.075 10.715 250.405 11.045 ;
        RECT 250.075 9.355 250.405 9.685 ;
        RECT 250.075 7.995 250.405 8.325 ;
        RECT 250.075 6.635 250.405 6.965 ;
        RECT 250.075 5.275 250.405 5.605 ;
        RECT 250.075 3.915 250.405 4.245 ;
        RECT 250.075 2.555 250.405 2.885 ;
        RECT 250.075 1.195 250.405 1.525 ;
        RECT 250.075 -0.165 250.405 0.165 ;
        RECT 250.08 -8.32 250.4 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 251.435 10.715 251.765 11.045 ;
        RECT 251.435 9.355 251.765 9.685 ;
        RECT 251.435 7.995 251.765 8.325 ;
        RECT 251.435 6.635 251.765 6.965 ;
        RECT 251.435 5.275 251.765 5.605 ;
        RECT 251.435 3.915 251.765 4.245 ;
        RECT 251.435 2.555 251.765 2.885 ;
        RECT 251.435 1.195 251.765 1.525 ;
        RECT 251.435 -0.165 251.765 0.165 ;
        RECT 251.44 -8.32 251.76 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.795 10.715 253.125 11.045 ;
        RECT 252.795 9.355 253.125 9.685 ;
        RECT 252.795 7.995 253.125 8.325 ;
        RECT 252.795 6.635 253.125 6.965 ;
        RECT 252.795 5.275 253.125 5.605 ;
        RECT 252.795 3.915 253.125 4.245 ;
        RECT 252.795 2.555 253.125 2.885 ;
        RECT 252.795 1.195 253.125 1.525 ;
        RECT 252.795 -0.165 253.125 0.165 ;
        RECT 252.8 -8.32 253.12 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 254.155 10.715 254.485 11.045 ;
        RECT 254.155 9.355 254.485 9.685 ;
        RECT 254.155 7.995 254.485 8.325 ;
        RECT 254.155 6.635 254.485 6.965 ;
        RECT 254.155 5.275 254.485 5.605 ;
        RECT 254.155 3.915 254.485 4.245 ;
        RECT 254.155 2.555 254.485 2.885 ;
        RECT 254.155 1.195 254.485 1.525 ;
        RECT 254.155 -0.165 254.485 0.165 ;
        RECT 254.16 -8.32 254.48 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 255.515 10.715 255.845 11.045 ;
        RECT 255.515 9.355 255.845 9.685 ;
        RECT 255.515 7.995 255.845 8.325 ;
        RECT 255.515 6.635 255.845 6.965 ;
        RECT 255.515 5.275 255.845 5.605 ;
        RECT 255.515 3.915 255.845 4.245 ;
        RECT 255.515 2.555 255.845 2.885 ;
        RECT 255.515 1.195 255.845 1.525 ;
        RECT 255.515 -0.165 255.845 0.165 ;
        RECT 255.52 -8.32 255.84 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 256.875 10.715 257.205 11.045 ;
        RECT 256.875 9.355 257.205 9.685 ;
        RECT 256.875 7.995 257.205 8.325 ;
        RECT 256.875 6.635 257.205 6.965 ;
        RECT 256.875 5.275 257.205 5.605 ;
        RECT 256.875 3.915 257.205 4.245 ;
        RECT 256.875 2.555 257.205 2.885 ;
        RECT 256.875 1.195 257.205 1.525 ;
        RECT 256.875 -0.165 257.205 0.165 ;
        RECT 256.88 -8.32 257.2 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.235 10.715 258.565 11.045 ;
        RECT 258.235 9.355 258.565 9.685 ;
        RECT 258.235 7.995 258.565 8.325 ;
        RECT 258.235 6.635 258.565 6.965 ;
        RECT 258.235 5.275 258.565 5.605 ;
        RECT 258.235 3.915 258.565 4.245 ;
        RECT 258.235 2.555 258.565 2.885 ;
        RECT 258.235 1.195 258.565 1.525 ;
        RECT 258.235 -0.165 258.565 0.165 ;
        RECT 258.24 -8.32 258.56 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 259.595 10.715 259.925 11.045 ;
        RECT 259.595 9.355 259.925 9.685 ;
        RECT 259.595 7.995 259.925 8.325 ;
        RECT 259.595 6.635 259.925 6.965 ;
        RECT 259.595 5.275 259.925 5.605 ;
        RECT 259.595 3.915 259.925 4.245 ;
        RECT 259.595 2.555 259.925 2.885 ;
        RECT 259.595 1.195 259.925 1.525 ;
        RECT 259.595 -0.165 259.925 0.165 ;
        RECT 259.6 -8.32 259.92 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.955 10.715 261.285 11.045 ;
        RECT 260.955 9.355 261.285 9.685 ;
        RECT 260.955 7.995 261.285 8.325 ;
        RECT 260.955 6.635 261.285 6.965 ;
        RECT 260.955 5.275 261.285 5.605 ;
        RECT 260.955 3.915 261.285 4.245 ;
        RECT 260.955 2.555 261.285 2.885 ;
        RECT 260.955 1.195 261.285 1.525 ;
        RECT 260.955 -0.165 261.285 0.165 ;
        RECT 260.96 -8.32 261.28 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.315 10.715 262.645 11.045 ;
        RECT 262.315 9.355 262.645 9.685 ;
        RECT 262.315 7.995 262.645 8.325 ;
        RECT 262.315 6.635 262.645 6.965 ;
        RECT 262.315 5.275 262.645 5.605 ;
        RECT 262.315 3.915 262.645 4.245 ;
        RECT 262.315 2.555 262.645 2.885 ;
        RECT 262.315 1.195 262.645 1.525 ;
        RECT 262.315 -0.165 262.645 0.165 ;
        RECT 262.32 -8.32 262.64 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 263.675 10.715 264.005 11.045 ;
        RECT 263.675 9.355 264.005 9.685 ;
        RECT 263.675 7.995 264.005 8.325 ;
        RECT 263.675 6.635 264.005 6.965 ;
        RECT 263.675 5.275 264.005 5.605 ;
        RECT 263.675 3.915 264.005 4.245 ;
        RECT 263.675 2.555 264.005 2.885 ;
        RECT 263.675 1.195 264.005 1.525 ;
        RECT 263.675 -0.165 264.005 0.165 ;
        RECT 263.68 -8.32 264 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 265.035 10.715 265.365 11.045 ;
        RECT 265.035 9.355 265.365 9.685 ;
        RECT 265.035 7.995 265.365 8.325 ;
        RECT 265.035 6.635 265.365 6.965 ;
        RECT 265.035 5.275 265.365 5.605 ;
        RECT 265.035 3.915 265.365 4.245 ;
        RECT 265.035 2.555 265.365 2.885 ;
        RECT 265.035 1.195 265.365 1.525 ;
        RECT 265.035 -0.165 265.365 0.165 ;
        RECT 265.04 -8.32 265.36 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 266.395 10.715 266.725 11.045 ;
        RECT 266.395 9.355 266.725 9.685 ;
        RECT 266.395 7.995 266.725 8.325 ;
        RECT 266.395 6.635 266.725 6.965 ;
        RECT 266.395 5.275 266.725 5.605 ;
        RECT 266.395 3.915 266.725 4.245 ;
        RECT 266.395 2.555 266.725 2.885 ;
        RECT 266.395 1.195 266.725 1.525 ;
        RECT 266.395 -0.165 266.725 0.165 ;
        RECT 266.4 -8.32 266.72 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 267.755 10.715 268.085 11.045 ;
        RECT 267.755 9.355 268.085 9.685 ;
        RECT 267.755 7.995 268.085 8.325 ;
        RECT 267.755 6.635 268.085 6.965 ;
        RECT 267.755 5.275 268.085 5.605 ;
        RECT 267.755 3.915 268.085 4.245 ;
        RECT 267.755 2.555 268.085 2.885 ;
        RECT 267.755 1.195 268.085 1.525 ;
        RECT 267.755 -0.165 268.085 0.165 ;
        RECT 267.76 -8.32 268.08 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.115 10.715 269.445 11.045 ;
        RECT 269.115 9.355 269.445 9.685 ;
        RECT 269.115 7.995 269.445 8.325 ;
        RECT 269.115 6.635 269.445 6.965 ;
        RECT 269.115 5.275 269.445 5.605 ;
        RECT 269.115 3.915 269.445 4.245 ;
        RECT 269.115 2.555 269.445 2.885 ;
        RECT 269.115 1.195 269.445 1.525 ;
        RECT 269.115 -0.165 269.445 0.165 ;
        RECT 269.12 -8.32 269.44 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 270.475 10.715 270.805 11.045 ;
        RECT 270.475 9.355 270.805 9.685 ;
        RECT 270.475 7.995 270.805 8.325 ;
        RECT 270.475 6.635 270.805 6.965 ;
        RECT 270.475 5.275 270.805 5.605 ;
        RECT 270.475 3.915 270.805 4.245 ;
        RECT 270.475 2.555 270.805 2.885 ;
        RECT 270.475 1.195 270.805 1.525 ;
        RECT 270.475 -0.165 270.805 0.165 ;
        RECT 270.48 -8.32 270.8 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.835 10.715 272.165 11.045 ;
        RECT 271.835 9.355 272.165 9.685 ;
        RECT 271.835 7.995 272.165 8.325 ;
        RECT 271.835 6.635 272.165 6.965 ;
        RECT 271.835 5.275 272.165 5.605 ;
        RECT 271.835 3.915 272.165 4.245 ;
        RECT 271.835 2.555 272.165 2.885 ;
        RECT 271.835 1.195 272.165 1.525 ;
        RECT 271.835 -0.165 272.165 0.165 ;
        RECT 271.84 -8.32 272.16 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.195 10.715 273.525 11.045 ;
        RECT 273.195 9.355 273.525 9.685 ;
        RECT 273.195 7.995 273.525 8.325 ;
        RECT 273.195 6.635 273.525 6.965 ;
        RECT 273.195 5.275 273.525 5.605 ;
        RECT 273.195 3.915 273.525 4.245 ;
        RECT 273.195 2.555 273.525 2.885 ;
        RECT 273.195 1.195 273.525 1.525 ;
        RECT 273.195 -0.165 273.525 0.165 ;
        RECT 273.2 -8.32 273.52 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 274.555 10.715 274.885 11.045 ;
        RECT 274.555 9.355 274.885 9.685 ;
        RECT 274.555 7.995 274.885 8.325 ;
        RECT 274.555 6.635 274.885 6.965 ;
        RECT 274.555 5.275 274.885 5.605 ;
        RECT 274.555 3.915 274.885 4.245 ;
        RECT 274.555 2.555 274.885 2.885 ;
        RECT 274.555 1.195 274.885 1.525 ;
        RECT 274.555 -0.165 274.885 0.165 ;
        RECT 274.56 -8.32 274.88 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.915 10.715 276.245 11.045 ;
        RECT 275.915 9.355 276.245 9.685 ;
        RECT 275.915 7.995 276.245 8.325 ;
        RECT 275.915 6.635 276.245 6.965 ;
        RECT 275.915 5.275 276.245 5.605 ;
        RECT 275.915 3.915 276.245 4.245 ;
        RECT 275.915 2.555 276.245 2.885 ;
        RECT 275.915 1.195 276.245 1.525 ;
        RECT 275.915 -0.165 276.245 0.165 ;
        RECT 275.92 -8.32 276.24 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 277.275 10.715 277.605 11.045 ;
        RECT 277.275 9.355 277.605 9.685 ;
        RECT 277.275 7.995 277.605 8.325 ;
        RECT 277.275 6.635 277.605 6.965 ;
        RECT 277.275 5.275 277.605 5.605 ;
        RECT 277.275 3.915 277.605 4.245 ;
        RECT 277.275 2.555 277.605 2.885 ;
        RECT 277.275 1.195 277.605 1.525 ;
        RECT 277.275 -0.165 277.605 0.165 ;
        RECT 277.28 -8.32 277.6 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 278.635 10.715 278.965 11.045 ;
        RECT 278.635 9.355 278.965 9.685 ;
        RECT 278.635 7.995 278.965 8.325 ;
        RECT 278.635 6.635 278.965 6.965 ;
        RECT 278.635 5.275 278.965 5.605 ;
        RECT 278.635 3.915 278.965 4.245 ;
        RECT 278.635 2.555 278.965 2.885 ;
        RECT 278.635 1.195 278.965 1.525 ;
        RECT 278.635 -0.165 278.965 0.165 ;
        RECT 278.64 -8.32 278.96 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.995 10.715 280.325 11.045 ;
        RECT 279.995 9.355 280.325 9.685 ;
        RECT 279.995 7.995 280.325 8.325 ;
        RECT 279.995 6.635 280.325 6.965 ;
        RECT 279.995 5.275 280.325 5.605 ;
        RECT 279.995 3.915 280.325 4.245 ;
        RECT 279.995 2.555 280.325 2.885 ;
        RECT 279.995 1.195 280.325 1.525 ;
        RECT 279.995 -0.165 280.325 0.165 ;
        RECT 280 -8.32 280.32 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 281.355 10.715 281.685 11.045 ;
        RECT 281.355 9.355 281.685 9.685 ;
        RECT 281.355 7.995 281.685 8.325 ;
        RECT 281.355 6.635 281.685 6.965 ;
        RECT 281.355 5.275 281.685 5.605 ;
        RECT 281.355 3.915 281.685 4.245 ;
        RECT 281.355 2.555 281.685 2.885 ;
        RECT 281.355 1.195 281.685 1.525 ;
        RECT 281.355 -0.165 281.685 0.165 ;
        RECT 281.36 -8.32 281.68 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.715 10.715 283.045 11.045 ;
        RECT 282.715 9.355 283.045 9.685 ;
        RECT 282.715 7.995 283.045 8.325 ;
        RECT 282.715 6.635 283.045 6.965 ;
        RECT 282.715 5.275 283.045 5.605 ;
        RECT 282.715 3.915 283.045 4.245 ;
        RECT 282.715 2.555 283.045 2.885 ;
        RECT 282.715 1.195 283.045 1.525 ;
        RECT 282.715 -0.165 283.045 0.165 ;
        RECT 282.72 -8.32 283.04 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 284.075 10.715 284.405 11.045 ;
        RECT 284.075 9.355 284.405 9.685 ;
        RECT 284.075 7.995 284.405 8.325 ;
        RECT 284.075 6.635 284.405 6.965 ;
        RECT 284.075 5.275 284.405 5.605 ;
        RECT 284.075 3.915 284.405 4.245 ;
        RECT 284.075 2.555 284.405 2.885 ;
        RECT 284.075 1.195 284.405 1.525 ;
        RECT 284.075 -0.165 284.405 0.165 ;
        RECT 284.08 -8.32 284.4 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 285.435 10.715 285.765 11.045 ;
        RECT 285.435 9.355 285.765 9.685 ;
        RECT 285.435 7.995 285.765 8.325 ;
        RECT 285.435 6.635 285.765 6.965 ;
        RECT 285.435 5.275 285.765 5.605 ;
        RECT 285.435 3.915 285.765 4.245 ;
        RECT 285.435 2.555 285.765 2.885 ;
        RECT 285.435 1.195 285.765 1.525 ;
        RECT 285.435 -0.165 285.765 0.165 ;
        RECT 285.44 -8.32 285.76 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.795 10.715 287.125 11.045 ;
        RECT 286.795 9.355 287.125 9.685 ;
        RECT 286.795 7.995 287.125 8.325 ;
        RECT 286.795 6.635 287.125 6.965 ;
        RECT 286.795 5.275 287.125 5.605 ;
        RECT 286.795 3.915 287.125 4.245 ;
        RECT 286.795 2.555 287.125 2.885 ;
        RECT 286.795 1.195 287.125 1.525 ;
        RECT 286.795 -0.165 287.125 0.165 ;
        RECT 286.8 -8.32 287.12 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.155 10.715 288.485 11.045 ;
        RECT 288.155 9.355 288.485 9.685 ;
        RECT 288.155 7.995 288.485 8.325 ;
        RECT 288.155 6.635 288.485 6.965 ;
        RECT 288.155 5.275 288.485 5.605 ;
        RECT 288.155 3.915 288.485 4.245 ;
        RECT 288.155 2.555 288.485 2.885 ;
        RECT 288.155 1.195 288.485 1.525 ;
        RECT 288.155 -0.165 288.485 0.165 ;
        RECT 288.16 -8.32 288.48 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 289.515 10.715 289.845 11.045 ;
        RECT 289.515 9.355 289.845 9.685 ;
        RECT 289.515 7.995 289.845 8.325 ;
        RECT 289.515 6.635 289.845 6.965 ;
        RECT 289.515 5.275 289.845 5.605 ;
        RECT 289.515 3.915 289.845 4.245 ;
        RECT 289.515 2.555 289.845 2.885 ;
        RECT 289.515 1.195 289.845 1.525 ;
        RECT 289.515 -0.165 289.845 0.165 ;
        RECT 289.52 -8.32 289.84 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.875 10.715 291.205 11.045 ;
        RECT 290.875 9.355 291.205 9.685 ;
        RECT 290.875 7.995 291.205 8.325 ;
        RECT 290.875 6.635 291.205 6.965 ;
        RECT 290.875 5.275 291.205 5.605 ;
        RECT 290.875 3.915 291.205 4.245 ;
        RECT 290.875 2.555 291.205 2.885 ;
        RECT 290.875 1.195 291.205 1.525 ;
        RECT 290.875 -0.165 291.205 0.165 ;
        RECT 290.88 -8.32 291.2 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.235 10.715 292.565 11.045 ;
        RECT 292.235 9.355 292.565 9.685 ;
        RECT 292.235 7.995 292.565 8.325 ;
        RECT 292.235 6.635 292.565 6.965 ;
        RECT 292.235 5.275 292.565 5.605 ;
        RECT 292.235 3.915 292.565 4.245 ;
        RECT 292.235 2.555 292.565 2.885 ;
        RECT 292.235 1.195 292.565 1.525 ;
        RECT 292.235 -0.165 292.565 0.165 ;
        RECT 292.24 -8.32 292.56 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 293.595 10.715 293.925 11.045 ;
        RECT 293.595 9.355 293.925 9.685 ;
        RECT 293.595 7.995 293.925 8.325 ;
        RECT 293.595 6.635 293.925 6.965 ;
        RECT 293.595 5.275 293.925 5.605 ;
        RECT 293.595 3.915 293.925 4.245 ;
        RECT 293.595 2.555 293.925 2.885 ;
        RECT 293.595 1.195 293.925 1.525 ;
        RECT 293.595 -0.165 293.925 0.165 ;
        RECT 293.6 -8.32 293.92 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.955 10.715 295.285 11.045 ;
        RECT 294.955 9.355 295.285 9.685 ;
        RECT 294.955 7.995 295.285 8.325 ;
        RECT 294.955 6.635 295.285 6.965 ;
        RECT 294.955 5.275 295.285 5.605 ;
        RECT 294.955 3.915 295.285 4.245 ;
        RECT 294.955 2.555 295.285 2.885 ;
        RECT 294.955 1.195 295.285 1.525 ;
        RECT 294.955 -0.165 295.285 0.165 ;
        RECT 294.96 -8.32 295.28 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 296.315 10.715 296.645 11.045 ;
        RECT 296.315 9.355 296.645 9.685 ;
        RECT 296.315 7.995 296.645 8.325 ;
        RECT 296.315 6.635 296.645 6.965 ;
        RECT 296.315 5.275 296.645 5.605 ;
        RECT 296.315 3.915 296.645 4.245 ;
        RECT 296.315 2.555 296.645 2.885 ;
        RECT 296.315 1.195 296.645 1.525 ;
        RECT 296.315 -0.165 296.645 0.165 ;
        RECT 296.32 -8.32 296.64 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 297.675 10.715 298.005 11.045 ;
        RECT 297.675 9.355 298.005 9.685 ;
        RECT 297.675 7.995 298.005 8.325 ;
        RECT 297.675 6.635 298.005 6.965 ;
        RECT 297.675 5.275 298.005 5.605 ;
        RECT 297.675 3.915 298.005 4.245 ;
        RECT 297.675 2.555 298.005 2.885 ;
        RECT 297.675 1.195 298.005 1.525 ;
        RECT 297.675 -0.165 298.005 0.165 ;
        RECT 297.68 -8.32 298 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 299.035 10.715 299.365 11.045 ;
        RECT 299.035 9.355 299.365 9.685 ;
        RECT 299.035 7.995 299.365 8.325 ;
        RECT 299.035 6.635 299.365 6.965 ;
        RECT 299.035 5.275 299.365 5.605 ;
        RECT 299.035 3.915 299.365 4.245 ;
        RECT 299.035 2.555 299.365 2.885 ;
        RECT 299.035 1.195 299.365 1.525 ;
        RECT 299.035 -0.165 299.365 0.165 ;
        RECT 299.04 -8.32 299.36 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 300.395 10.715 300.725 11.045 ;
        RECT 300.395 9.355 300.725 9.685 ;
        RECT 300.395 7.995 300.725 8.325 ;
        RECT 300.395 6.635 300.725 6.965 ;
        RECT 300.395 5.275 300.725 5.605 ;
        RECT 300.395 3.915 300.725 4.245 ;
        RECT 300.395 2.555 300.725 2.885 ;
        RECT 300.395 1.195 300.725 1.525 ;
        RECT 300.395 -0.165 300.725 0.165 ;
        RECT 300.4 -8.32 300.72 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.755 10.715 302.085 11.045 ;
        RECT 301.755 9.355 302.085 9.685 ;
        RECT 301.755 7.995 302.085 8.325 ;
        RECT 301.755 6.635 302.085 6.965 ;
        RECT 301.755 5.275 302.085 5.605 ;
        RECT 301.755 3.915 302.085 4.245 ;
        RECT 301.755 2.555 302.085 2.885 ;
        RECT 301.755 1.195 302.085 1.525 ;
        RECT 301.755 -0.165 302.085 0.165 ;
        RECT 301.76 -8.32 302.08 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.115 10.715 303.445 11.045 ;
        RECT 303.115 9.355 303.445 9.685 ;
        RECT 303.115 7.995 303.445 8.325 ;
        RECT 303.115 6.635 303.445 6.965 ;
        RECT 303.115 5.275 303.445 5.605 ;
        RECT 303.115 3.915 303.445 4.245 ;
        RECT 303.115 2.555 303.445 2.885 ;
        RECT 303.115 1.195 303.445 1.525 ;
        RECT 303.115 -0.165 303.445 0.165 ;
        RECT 303.12 -8.32 303.44 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 304.475 10.715 304.805 11.045 ;
        RECT 304.475 9.355 304.805 9.685 ;
        RECT 304.475 7.995 304.805 8.325 ;
        RECT 304.475 6.635 304.805 6.965 ;
        RECT 304.475 5.275 304.805 5.605 ;
        RECT 304.475 3.915 304.805 4.245 ;
        RECT 304.475 2.555 304.805 2.885 ;
        RECT 304.475 1.195 304.805 1.525 ;
        RECT 304.475 -0.165 304.805 0.165 ;
        RECT 304.48 -8.32 304.8 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.835 10.715 306.165 11.045 ;
        RECT 305.835 9.355 306.165 9.685 ;
        RECT 305.835 7.995 306.165 8.325 ;
        RECT 305.835 6.635 306.165 6.965 ;
        RECT 305.835 5.275 306.165 5.605 ;
        RECT 305.835 3.915 306.165 4.245 ;
        RECT 305.835 2.555 306.165 2.885 ;
        RECT 305.835 1.195 306.165 1.525 ;
        RECT 305.835 -0.165 306.165 0.165 ;
        RECT 305.84 -8.32 306.16 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.195 10.715 307.525 11.045 ;
        RECT 307.195 9.355 307.525 9.685 ;
        RECT 307.195 7.995 307.525 8.325 ;
        RECT 307.195 6.635 307.525 6.965 ;
        RECT 307.195 5.275 307.525 5.605 ;
        RECT 307.195 3.915 307.525 4.245 ;
        RECT 307.195 2.555 307.525 2.885 ;
        RECT 307.195 1.195 307.525 1.525 ;
        RECT 307.195 -0.165 307.525 0.165 ;
        RECT 307.2 -8.32 307.52 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 308.555 10.715 308.885 11.045 ;
        RECT 308.555 9.355 308.885 9.685 ;
        RECT 308.555 7.995 308.885 8.325 ;
        RECT 308.555 6.635 308.885 6.965 ;
        RECT 308.555 5.275 308.885 5.605 ;
        RECT 308.555 3.915 308.885 4.245 ;
        RECT 308.555 2.555 308.885 2.885 ;
        RECT 308.555 1.195 308.885 1.525 ;
        RECT 308.555 -0.165 308.885 0.165 ;
        RECT 308.56 -8.32 308.88 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.915 10.715 310.245 11.045 ;
        RECT 309.915 9.355 310.245 9.685 ;
        RECT 309.915 7.995 310.245 8.325 ;
        RECT 309.915 6.635 310.245 6.965 ;
        RECT 309.915 5.275 310.245 5.605 ;
        RECT 309.915 3.915 310.245 4.245 ;
        RECT 309.915 2.555 310.245 2.885 ;
        RECT 309.915 1.195 310.245 1.525 ;
        RECT 309.915 -0.165 310.245 0.165 ;
        RECT 309.92 -8.32 310.24 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 311.275 10.715 311.605 11.045 ;
        RECT 311.275 9.355 311.605 9.685 ;
        RECT 311.275 7.995 311.605 8.325 ;
        RECT 311.275 6.635 311.605 6.965 ;
        RECT 311.275 5.275 311.605 5.605 ;
        RECT 311.275 3.915 311.605 4.245 ;
        RECT 311.275 2.555 311.605 2.885 ;
        RECT 311.275 1.195 311.605 1.525 ;
        RECT 311.275 -0.165 311.605 0.165 ;
        RECT 311.28 -8.32 311.6 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 312.635 10.715 312.965 11.045 ;
        RECT 312.635 9.355 312.965 9.685 ;
        RECT 312.635 7.995 312.965 8.325 ;
        RECT 312.635 6.635 312.965 6.965 ;
        RECT 312.635 5.275 312.965 5.605 ;
        RECT 312.635 3.915 312.965 4.245 ;
        RECT 312.635 2.555 312.965 2.885 ;
        RECT 312.635 1.195 312.965 1.525 ;
        RECT 312.635 -0.165 312.965 0.165 ;
        RECT 312.64 -8.32 312.96 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.995 10.715 314.325 11.045 ;
        RECT 313.995 9.355 314.325 9.685 ;
        RECT 313.995 7.995 314.325 8.325 ;
        RECT 313.995 6.635 314.325 6.965 ;
        RECT 313.995 5.275 314.325 5.605 ;
        RECT 313.995 3.915 314.325 4.245 ;
        RECT 313.995 2.555 314.325 2.885 ;
        RECT 313.995 1.195 314.325 1.525 ;
        RECT 313.995 -0.165 314.325 0.165 ;
        RECT 314 -8.32 314.32 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 315.355 10.715 315.685 11.045 ;
        RECT 315.355 9.355 315.685 9.685 ;
        RECT 315.355 7.995 315.685 8.325 ;
        RECT 315.355 6.635 315.685 6.965 ;
        RECT 315.355 5.275 315.685 5.605 ;
        RECT 315.355 3.915 315.685 4.245 ;
        RECT 315.355 2.555 315.685 2.885 ;
        RECT 315.355 1.195 315.685 1.525 ;
        RECT 315.355 -0.165 315.685 0.165 ;
        RECT 315.36 -8.32 315.68 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 316.715 10.715 317.045 11.045 ;
        RECT 316.715 9.355 317.045 9.685 ;
        RECT 316.715 7.995 317.045 8.325 ;
        RECT 316.715 6.635 317.045 6.965 ;
        RECT 316.715 5.275 317.045 5.605 ;
        RECT 316.715 3.915 317.045 4.245 ;
        RECT 316.715 2.555 317.045 2.885 ;
        RECT 316.715 1.195 317.045 1.525 ;
        RECT 316.715 -0.165 317.045 0.165 ;
        RECT 316.72 -8.32 317.04 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.075 10.715 318.405 11.045 ;
        RECT 318.075 9.355 318.405 9.685 ;
        RECT 318.075 7.995 318.405 8.325 ;
        RECT 318.075 6.635 318.405 6.965 ;
        RECT 318.075 5.275 318.405 5.605 ;
        RECT 318.075 3.915 318.405 4.245 ;
        RECT 318.075 2.555 318.405 2.885 ;
        RECT 318.075 1.195 318.405 1.525 ;
        RECT 318.075 -0.165 318.405 0.165 ;
        RECT 318.08 -8.32 318.4 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 319.435 10.715 319.765 11.045 ;
        RECT 319.435 9.355 319.765 9.685 ;
        RECT 319.435 7.995 319.765 8.325 ;
        RECT 319.435 6.635 319.765 6.965 ;
        RECT 319.435 5.275 319.765 5.605 ;
        RECT 319.435 3.915 319.765 4.245 ;
        RECT 319.435 2.555 319.765 2.885 ;
        RECT 319.435 1.195 319.765 1.525 ;
        RECT 319.435 -0.165 319.765 0.165 ;
        RECT 319.44 -8.32 319.76 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 320.795 10.715 321.125 11.045 ;
        RECT 320.795 9.355 321.125 9.685 ;
        RECT 320.795 7.995 321.125 8.325 ;
        RECT 320.795 6.635 321.125 6.965 ;
        RECT 320.795 5.275 321.125 5.605 ;
        RECT 320.795 3.915 321.125 4.245 ;
        RECT 320.795 2.555 321.125 2.885 ;
        RECT 320.795 1.195 321.125 1.525 ;
        RECT 320.795 -0.165 321.125 0.165 ;
        RECT 320.8 -8.32 321.12 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 322.155 10.715 322.485 11.045 ;
        RECT 322.155 9.355 322.485 9.685 ;
        RECT 322.155 7.995 322.485 8.325 ;
        RECT 322.155 6.635 322.485 6.965 ;
        RECT 322.155 5.275 322.485 5.605 ;
        RECT 322.155 3.915 322.485 4.245 ;
        RECT 322.155 2.555 322.485 2.885 ;
        RECT 322.155 1.195 322.485 1.525 ;
        RECT 322.155 -0.165 322.485 0.165 ;
        RECT 322.16 -8.32 322.48 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 323.515 10.715 323.845 11.045 ;
        RECT 323.515 9.355 323.845 9.685 ;
        RECT 323.515 7.995 323.845 8.325 ;
        RECT 323.515 6.635 323.845 6.965 ;
        RECT 323.515 5.275 323.845 5.605 ;
        RECT 323.515 3.915 323.845 4.245 ;
        RECT 323.515 2.555 323.845 2.885 ;
        RECT 323.515 1.195 323.845 1.525 ;
        RECT 323.515 -0.165 323.845 0.165 ;
        RECT 323.52 -8.32 323.84 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.875 10.715 325.205 11.045 ;
        RECT 324.875 9.355 325.205 9.685 ;
        RECT 324.875 7.995 325.205 8.325 ;
        RECT 324.875 6.635 325.205 6.965 ;
        RECT 324.875 5.275 325.205 5.605 ;
        RECT 324.875 3.915 325.205 4.245 ;
        RECT 324.875 2.555 325.205 2.885 ;
        RECT 324.875 1.195 325.205 1.525 ;
        RECT 324.875 -0.165 325.205 0.165 ;
        RECT 324.88 -8.32 325.2 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 326.235 10.715 326.565 11.045 ;
        RECT 326.235 9.355 326.565 9.685 ;
        RECT 326.235 7.995 326.565 8.325 ;
        RECT 326.235 6.635 326.565 6.965 ;
        RECT 326.235 5.275 326.565 5.605 ;
        RECT 326.235 3.915 326.565 4.245 ;
        RECT 326.235 2.555 326.565 2.885 ;
        RECT 326.235 1.195 326.565 1.525 ;
        RECT 326.235 -0.165 326.565 0.165 ;
        RECT 326.24 -8.32 326.56 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 327.595 10.715 327.925 11.045 ;
        RECT 327.595 9.355 327.925 9.685 ;
        RECT 327.595 7.995 327.925 8.325 ;
        RECT 327.595 6.635 327.925 6.965 ;
        RECT 327.595 5.275 327.925 5.605 ;
        RECT 327.595 3.915 327.925 4.245 ;
        RECT 327.595 2.555 327.925 2.885 ;
        RECT 327.595 1.195 327.925 1.525 ;
        RECT 327.595 -0.165 327.925 0.165 ;
        RECT 327.6 -8.32 327.92 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 328.955 10.715 329.285 11.045 ;
        RECT 328.955 9.355 329.285 9.685 ;
        RECT 328.955 7.995 329.285 8.325 ;
        RECT 328.955 6.635 329.285 6.965 ;
        RECT 328.955 5.275 329.285 5.605 ;
        RECT 328.955 3.915 329.285 4.245 ;
        RECT 328.955 2.555 329.285 2.885 ;
        RECT 328.955 1.195 329.285 1.525 ;
        RECT 328.955 -0.165 329.285 0.165 ;
        RECT 328.96 -8.32 329.28 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.315 10.715 330.645 11.045 ;
        RECT 330.315 9.355 330.645 9.685 ;
        RECT 330.315 7.995 330.645 8.325 ;
        RECT 330.315 6.635 330.645 6.965 ;
        RECT 330.315 5.275 330.645 5.605 ;
        RECT 330.315 3.915 330.645 4.245 ;
        RECT 330.315 2.555 330.645 2.885 ;
        RECT 330.315 1.195 330.645 1.525 ;
        RECT 330.315 -0.165 330.645 0.165 ;
        RECT 330.32 -8.32 330.64 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 331.675 10.715 332.005 11.045 ;
        RECT 331.675 9.355 332.005 9.685 ;
        RECT 331.675 7.995 332.005 8.325 ;
        RECT 331.675 6.635 332.005 6.965 ;
        RECT 331.675 5.275 332.005 5.605 ;
        RECT 331.675 3.915 332.005 4.245 ;
        RECT 331.675 2.555 332.005 2.885 ;
        RECT 331.675 1.195 332.005 1.525 ;
        RECT 331.675 -0.165 332.005 0.165 ;
        RECT 331.68 -8.32 332 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 333.035 10.715 333.365 11.045 ;
        RECT 333.035 9.355 333.365 9.685 ;
        RECT 333.035 7.995 333.365 8.325 ;
        RECT 333.035 6.635 333.365 6.965 ;
        RECT 333.035 5.275 333.365 5.605 ;
        RECT 333.035 3.915 333.365 4.245 ;
        RECT 333.035 2.555 333.365 2.885 ;
        RECT 333.035 1.195 333.365 1.525 ;
        RECT 333.035 -0.165 333.365 0.165 ;
        RECT 333.04 -8.32 333.36 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 334.395 10.715 334.725 11.045 ;
        RECT 334.395 9.355 334.725 9.685 ;
        RECT 334.395 7.995 334.725 8.325 ;
        RECT 334.395 6.635 334.725 6.965 ;
        RECT 334.395 5.275 334.725 5.605 ;
        RECT 334.395 3.915 334.725 4.245 ;
        RECT 334.395 2.555 334.725 2.885 ;
        RECT 334.395 1.195 334.725 1.525 ;
        RECT 334.395 -0.165 334.725 0.165 ;
        RECT 334.4 -8.32 334.72 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.755 10.715 336.085 11.045 ;
        RECT 335.755 9.355 336.085 9.685 ;
        RECT 335.755 7.995 336.085 8.325 ;
        RECT 335.755 6.635 336.085 6.965 ;
        RECT 335.755 5.275 336.085 5.605 ;
        RECT 335.755 3.915 336.085 4.245 ;
        RECT 335.755 2.555 336.085 2.885 ;
        RECT 335.755 1.195 336.085 1.525 ;
        RECT 335.755 -0.165 336.085 0.165 ;
        RECT 335.76 -8.32 336.08 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 337.115 10.715 337.445 11.045 ;
        RECT 337.115 9.355 337.445 9.685 ;
        RECT 337.115 7.995 337.445 8.325 ;
        RECT 337.115 6.635 337.445 6.965 ;
        RECT 337.115 5.275 337.445 5.605 ;
        RECT 337.115 3.915 337.445 4.245 ;
        RECT 337.115 2.555 337.445 2.885 ;
        RECT 337.115 1.195 337.445 1.525 ;
        RECT 337.115 -0.165 337.445 0.165 ;
        RECT 337.12 -8.32 337.44 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 338.475 10.715 338.805 11.045 ;
        RECT 338.475 9.355 338.805 9.685 ;
        RECT 338.475 7.995 338.805 8.325 ;
        RECT 338.475 6.635 338.805 6.965 ;
        RECT 338.475 5.275 338.805 5.605 ;
        RECT 338.475 3.915 338.805 4.245 ;
        RECT 338.475 2.555 338.805 2.885 ;
        RECT 338.475 1.195 338.805 1.525 ;
        RECT 338.475 -0.165 338.805 0.165 ;
        RECT 338.48 -8.32 338.8 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 339.835 10.715 340.165 11.045 ;
        RECT 339.835 9.355 340.165 9.685 ;
        RECT 339.835 7.995 340.165 8.325 ;
        RECT 339.835 6.635 340.165 6.965 ;
        RECT 339.835 5.275 340.165 5.605 ;
        RECT 339.835 3.915 340.165 4.245 ;
        RECT 339.835 2.555 340.165 2.885 ;
        RECT 339.835 1.195 340.165 1.525 ;
        RECT 339.835 -0.165 340.165 0.165 ;
        RECT 339.84 -8.32 340.16 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 341.195 10.715 341.525 11.045 ;
        RECT 341.195 9.355 341.525 9.685 ;
        RECT 341.195 7.995 341.525 8.325 ;
        RECT 341.195 6.635 341.525 6.965 ;
        RECT 341.195 5.275 341.525 5.605 ;
        RECT 341.195 3.915 341.525 4.245 ;
        RECT 341.195 2.555 341.525 2.885 ;
        RECT 341.195 1.195 341.525 1.525 ;
        RECT 341.195 -0.165 341.525 0.165 ;
        RECT 341.2 -8.32 341.52 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 342.555 10.715 342.885 11.045 ;
        RECT 342.555 9.355 342.885 9.685 ;
        RECT 342.555 7.995 342.885 8.325 ;
        RECT 342.555 6.635 342.885 6.965 ;
        RECT 342.555 5.275 342.885 5.605 ;
        RECT 342.555 3.915 342.885 4.245 ;
        RECT 342.555 2.555 342.885 2.885 ;
        RECT 342.555 1.195 342.885 1.525 ;
        RECT 342.555 -0.165 342.885 0.165 ;
        RECT 342.56 -8.32 342.88 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 343.915 10.715 344.245 11.045 ;
        RECT 343.915 9.355 344.245 9.685 ;
        RECT 343.915 7.995 344.245 8.325 ;
        RECT 343.915 6.635 344.245 6.965 ;
        RECT 343.915 5.275 344.245 5.605 ;
        RECT 343.915 3.915 344.245 4.245 ;
        RECT 343.915 2.555 344.245 2.885 ;
        RECT 343.915 1.195 344.245 1.525 ;
        RECT 343.915 -0.165 344.245 0.165 ;
        RECT 343.92 -8.32 344.24 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 345.275 10.715 345.605 11.045 ;
        RECT 345.275 9.355 345.605 9.685 ;
        RECT 345.275 7.995 345.605 8.325 ;
        RECT 345.275 6.635 345.605 6.965 ;
        RECT 345.275 5.275 345.605 5.605 ;
        RECT 345.275 3.915 345.605 4.245 ;
        RECT 345.275 2.555 345.605 2.885 ;
        RECT 345.275 1.195 345.605 1.525 ;
        RECT 345.275 -0.165 345.605 0.165 ;
        RECT 345.28 -8.32 345.6 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 346.635 10.715 346.965 11.045 ;
        RECT 346.635 9.355 346.965 9.685 ;
        RECT 346.635 7.995 346.965 8.325 ;
        RECT 346.635 6.635 346.965 6.965 ;
        RECT 346.635 5.275 346.965 5.605 ;
        RECT 346.635 3.915 346.965 4.245 ;
        RECT 346.635 2.555 346.965 2.885 ;
        RECT 346.635 1.195 346.965 1.525 ;
        RECT 346.635 -0.165 346.965 0.165 ;
        RECT 346.64 -8.32 346.96 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 347.995 10.715 348.325 11.045 ;
        RECT 347.995 9.355 348.325 9.685 ;
        RECT 347.995 7.995 348.325 8.325 ;
        RECT 347.995 6.635 348.325 6.965 ;
        RECT 347.995 5.275 348.325 5.605 ;
        RECT 347.995 3.915 348.325 4.245 ;
        RECT 347.995 2.555 348.325 2.885 ;
        RECT 347.995 1.195 348.325 1.525 ;
        RECT 347.995 -0.165 348.325 0.165 ;
        RECT 348 -8.32 348.32 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 349.355 10.715 349.685 11.045 ;
        RECT 349.355 9.355 349.685 9.685 ;
        RECT 349.355 7.995 349.685 8.325 ;
        RECT 349.355 6.635 349.685 6.965 ;
        RECT 349.355 5.275 349.685 5.605 ;
        RECT 349.355 3.915 349.685 4.245 ;
        RECT 349.355 2.555 349.685 2.885 ;
        RECT 349.355 1.195 349.685 1.525 ;
        RECT 349.355 -0.165 349.685 0.165 ;
        RECT 349.36 -8.32 349.68 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 350.715 10.715 351.045 11.045 ;
        RECT 350.715 9.355 351.045 9.685 ;
        RECT 350.715 7.995 351.045 8.325 ;
        RECT 350.715 6.635 351.045 6.965 ;
        RECT 350.715 5.275 351.045 5.605 ;
        RECT 350.715 3.915 351.045 4.245 ;
        RECT 350.715 2.555 351.045 2.885 ;
        RECT 350.715 1.195 351.045 1.525 ;
        RECT 350.715 -0.165 351.045 0.165 ;
        RECT 350.72 -8.32 351.04 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 352.075 10.715 352.405 11.045 ;
        RECT 352.075 9.355 352.405 9.685 ;
        RECT 352.075 7.995 352.405 8.325 ;
        RECT 352.075 6.635 352.405 6.965 ;
        RECT 352.075 5.275 352.405 5.605 ;
        RECT 352.075 3.915 352.405 4.245 ;
        RECT 352.075 2.555 352.405 2.885 ;
        RECT 352.075 1.195 352.405 1.525 ;
        RECT 352.075 -0.165 352.405 0.165 ;
        RECT 352.08 -8.32 352.4 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 353.435 10.715 353.765 11.045 ;
        RECT 353.435 9.355 353.765 9.685 ;
        RECT 353.435 7.995 353.765 8.325 ;
        RECT 353.435 6.635 353.765 6.965 ;
        RECT 353.435 5.275 353.765 5.605 ;
        RECT 353.435 3.915 353.765 4.245 ;
        RECT 353.435 2.555 353.765 2.885 ;
        RECT 353.435 1.195 353.765 1.525 ;
        RECT 353.435 -0.165 353.765 0.165 ;
        RECT 353.44 -8.32 353.76 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.795 10.715 355.125 11.045 ;
        RECT 354.795 9.355 355.125 9.685 ;
        RECT 354.795 7.995 355.125 8.325 ;
        RECT 354.795 6.635 355.125 6.965 ;
        RECT 354.795 5.275 355.125 5.605 ;
        RECT 354.795 3.915 355.125 4.245 ;
        RECT 354.795 2.555 355.125 2.885 ;
        RECT 354.795 1.195 355.125 1.525 ;
        RECT 354.795 -0.165 355.125 0.165 ;
        RECT 354.8 -8.32 355.12 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 356.155 10.715 356.485 11.045 ;
        RECT 356.155 9.355 356.485 9.685 ;
        RECT 356.155 7.995 356.485 8.325 ;
        RECT 356.155 6.635 356.485 6.965 ;
        RECT 356.155 5.275 356.485 5.605 ;
        RECT 356.155 3.915 356.485 4.245 ;
        RECT 356.155 2.555 356.485 2.885 ;
        RECT 356.155 1.195 356.485 1.525 ;
        RECT 356.155 -0.165 356.485 0.165 ;
        RECT 356.16 -8.32 356.48 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 357.515 10.715 357.845 11.045 ;
        RECT 357.515 9.355 357.845 9.685 ;
        RECT 357.515 7.995 357.845 8.325 ;
        RECT 357.515 6.635 357.845 6.965 ;
        RECT 357.515 5.275 357.845 5.605 ;
        RECT 357.515 3.915 357.845 4.245 ;
        RECT 357.515 2.555 357.845 2.885 ;
        RECT 357.515 1.195 357.845 1.525 ;
        RECT 357.515 -0.165 357.845 0.165 ;
        RECT 357.52 -8.32 357.84 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 358.875 10.715 359.205 11.045 ;
        RECT 358.875 9.355 359.205 9.685 ;
        RECT 358.875 7.995 359.205 8.325 ;
        RECT 358.875 6.635 359.205 6.965 ;
        RECT 358.875 5.275 359.205 5.605 ;
        RECT 358.875 3.915 359.205 4.245 ;
        RECT 358.875 2.555 359.205 2.885 ;
        RECT 358.875 1.195 359.205 1.525 ;
        RECT 358.875 -0.165 359.205 0.165 ;
        RECT 358.88 -8.32 359.2 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 360.235 10.715 360.565 11.045 ;
        RECT 360.235 9.355 360.565 9.685 ;
        RECT 360.235 7.995 360.565 8.325 ;
        RECT 360.235 6.635 360.565 6.965 ;
        RECT 360.235 5.275 360.565 5.605 ;
        RECT 360.235 3.915 360.565 4.245 ;
        RECT 360.235 2.555 360.565 2.885 ;
        RECT 360.235 1.195 360.565 1.525 ;
        RECT 360.235 -0.165 360.565 0.165 ;
        RECT 360.24 -8.32 360.56 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 361.595 9.355 361.925 9.685 ;
        RECT 361.595 7.995 361.925 8.325 ;
        RECT 361.595 6.635 361.925 6.965 ;
        RECT 361.595 5.275 361.925 5.605 ;
        RECT 361.595 3.915 361.925 4.245 ;
        RECT 361.595 2.555 361.925 2.885 ;
        RECT 361.595 1.195 361.925 1.525 ;
        RECT 361.595 -0.165 361.925 0.165 ;
        RECT 361.6 -8.32 361.92 15.8 ;
        RECT 361.595 10.715 361.925 11.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.955 10.715 91.285 11.045 ;
        RECT 90.955 9.355 91.285 9.685 ;
        RECT 90.955 7.995 91.285 8.325 ;
        RECT 90.955 6.635 91.285 6.965 ;
        RECT 90.955 5.275 91.285 5.605 ;
        RECT 90.955 3.915 91.285 4.245 ;
        RECT 90.955 2.555 91.285 2.885 ;
        RECT 90.955 1.195 91.285 1.525 ;
        RECT 90.955 -0.165 91.285 0.165 ;
        RECT 90.96 -8.32 91.28 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.315 10.715 92.645 11.045 ;
        RECT 92.315 9.355 92.645 9.685 ;
        RECT 92.315 7.995 92.645 8.325 ;
        RECT 92.315 6.635 92.645 6.965 ;
        RECT 92.315 5.275 92.645 5.605 ;
        RECT 92.315 3.915 92.645 4.245 ;
        RECT 92.315 2.555 92.645 2.885 ;
        RECT 92.315 1.195 92.645 1.525 ;
        RECT 92.315 -0.165 92.645 0.165 ;
        RECT 92.32 -8.32 92.64 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.675 10.715 94.005 11.045 ;
        RECT 93.675 9.355 94.005 9.685 ;
        RECT 93.675 7.995 94.005 8.325 ;
        RECT 93.675 6.635 94.005 6.965 ;
        RECT 93.675 5.275 94.005 5.605 ;
        RECT 93.675 3.915 94.005 4.245 ;
        RECT 93.675 2.555 94.005 2.885 ;
        RECT 93.675 1.195 94.005 1.525 ;
        RECT 93.675 -0.165 94.005 0.165 ;
        RECT 93.68 -8.32 94 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.035 10.715 95.365 11.045 ;
        RECT 95.035 9.355 95.365 9.685 ;
        RECT 95.035 7.995 95.365 8.325 ;
        RECT 95.035 6.635 95.365 6.965 ;
        RECT 95.035 5.275 95.365 5.605 ;
        RECT 95.035 3.915 95.365 4.245 ;
        RECT 95.035 2.555 95.365 2.885 ;
        RECT 95.035 1.195 95.365 1.525 ;
        RECT 95.035 -0.165 95.365 0.165 ;
        RECT 95.04 -8.32 95.36 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.395 10.715 96.725 11.045 ;
        RECT 96.395 9.355 96.725 9.685 ;
        RECT 96.395 7.995 96.725 8.325 ;
        RECT 96.395 6.635 96.725 6.965 ;
        RECT 96.395 5.275 96.725 5.605 ;
        RECT 96.395 3.915 96.725 4.245 ;
        RECT 96.395 2.555 96.725 2.885 ;
        RECT 96.395 1.195 96.725 1.525 ;
        RECT 96.395 -0.165 96.725 0.165 ;
        RECT 96.4 -8.32 96.72 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.755 10.715 98.085 11.045 ;
        RECT 97.755 9.355 98.085 9.685 ;
        RECT 97.755 7.995 98.085 8.325 ;
        RECT 97.755 6.635 98.085 6.965 ;
        RECT 97.755 5.275 98.085 5.605 ;
        RECT 97.755 3.915 98.085 4.245 ;
        RECT 97.755 2.555 98.085 2.885 ;
        RECT 97.755 1.195 98.085 1.525 ;
        RECT 97.755 -0.165 98.085 0.165 ;
        RECT 97.76 -8.32 98.08 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.115 10.715 99.445 11.045 ;
        RECT 99.115 9.355 99.445 9.685 ;
        RECT 99.115 7.995 99.445 8.325 ;
        RECT 99.115 6.635 99.445 6.965 ;
        RECT 99.115 5.275 99.445 5.605 ;
        RECT 99.115 3.915 99.445 4.245 ;
        RECT 99.115 2.555 99.445 2.885 ;
        RECT 99.115 1.195 99.445 1.525 ;
        RECT 99.115 -0.165 99.445 0.165 ;
        RECT 99.12 -8.32 99.44 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.475 10.715 100.805 11.045 ;
        RECT 100.475 9.355 100.805 9.685 ;
        RECT 100.475 7.995 100.805 8.325 ;
        RECT 100.475 6.635 100.805 6.965 ;
        RECT 100.475 5.275 100.805 5.605 ;
        RECT 100.475 3.915 100.805 4.245 ;
        RECT 100.475 2.555 100.805 2.885 ;
        RECT 100.475 1.195 100.805 1.525 ;
        RECT 100.475 -0.165 100.805 0.165 ;
        RECT 100.48 -8.32 100.8 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.835 10.715 102.165 11.045 ;
        RECT 101.835 9.355 102.165 9.685 ;
        RECT 101.835 7.995 102.165 8.325 ;
        RECT 101.835 6.635 102.165 6.965 ;
        RECT 101.835 5.275 102.165 5.605 ;
        RECT 101.835 3.915 102.165 4.245 ;
        RECT 101.835 2.555 102.165 2.885 ;
        RECT 101.835 1.195 102.165 1.525 ;
        RECT 101.835 -0.165 102.165 0.165 ;
        RECT 101.84 -8.32 102.16 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.195 10.715 103.525 11.045 ;
        RECT 103.195 9.355 103.525 9.685 ;
        RECT 103.195 7.995 103.525 8.325 ;
        RECT 103.195 6.635 103.525 6.965 ;
        RECT 103.195 5.275 103.525 5.605 ;
        RECT 103.195 3.915 103.525 4.245 ;
        RECT 103.195 2.555 103.525 2.885 ;
        RECT 103.195 1.195 103.525 1.525 ;
        RECT 103.195 -0.165 103.525 0.165 ;
        RECT 103.2 -8.32 103.52 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 104.555 10.715 104.885 11.045 ;
        RECT 104.555 9.355 104.885 9.685 ;
        RECT 104.555 7.995 104.885 8.325 ;
        RECT 104.555 6.635 104.885 6.965 ;
        RECT 104.555 5.275 104.885 5.605 ;
        RECT 104.555 3.915 104.885 4.245 ;
        RECT 104.555 2.555 104.885 2.885 ;
        RECT 104.555 1.195 104.885 1.525 ;
        RECT 104.555 -0.165 104.885 0.165 ;
        RECT 104.56 -8.32 104.88 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.915 10.715 106.245 11.045 ;
        RECT 105.915 9.355 106.245 9.685 ;
        RECT 105.915 7.995 106.245 8.325 ;
        RECT 105.915 6.635 106.245 6.965 ;
        RECT 105.915 5.275 106.245 5.605 ;
        RECT 105.915 3.915 106.245 4.245 ;
        RECT 105.915 2.555 106.245 2.885 ;
        RECT 105.915 1.195 106.245 1.525 ;
        RECT 105.915 -0.165 106.245 0.165 ;
        RECT 105.92 -8.32 106.24 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.275 10.715 107.605 11.045 ;
        RECT 107.275 9.355 107.605 9.685 ;
        RECT 107.275 7.995 107.605 8.325 ;
        RECT 107.275 6.635 107.605 6.965 ;
        RECT 107.275 5.275 107.605 5.605 ;
        RECT 107.275 3.915 107.605 4.245 ;
        RECT 107.275 2.555 107.605 2.885 ;
        RECT 107.275 1.195 107.605 1.525 ;
        RECT 107.275 -0.165 107.605 0.165 ;
        RECT 107.28 -8.32 107.6 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.635 10.715 108.965 11.045 ;
        RECT 108.635 9.355 108.965 9.685 ;
        RECT 108.635 7.995 108.965 8.325 ;
        RECT 108.635 6.635 108.965 6.965 ;
        RECT 108.635 5.275 108.965 5.605 ;
        RECT 108.635 3.915 108.965 4.245 ;
        RECT 108.635 2.555 108.965 2.885 ;
        RECT 108.635 1.195 108.965 1.525 ;
        RECT 108.635 -0.165 108.965 0.165 ;
        RECT 108.64 -8.32 108.96 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.995 10.715 110.325 11.045 ;
        RECT 109.995 9.355 110.325 9.685 ;
        RECT 109.995 7.995 110.325 8.325 ;
        RECT 109.995 6.635 110.325 6.965 ;
        RECT 109.995 5.275 110.325 5.605 ;
        RECT 109.995 3.915 110.325 4.245 ;
        RECT 109.995 2.555 110.325 2.885 ;
        RECT 109.995 1.195 110.325 1.525 ;
        RECT 109.995 -0.165 110.325 0.165 ;
        RECT 110 -8.32 110.32 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.355 10.715 111.685 11.045 ;
        RECT 111.355 9.355 111.685 9.685 ;
        RECT 111.355 7.995 111.685 8.325 ;
        RECT 111.355 6.635 111.685 6.965 ;
        RECT 111.355 5.275 111.685 5.605 ;
        RECT 111.355 3.915 111.685 4.245 ;
        RECT 111.355 2.555 111.685 2.885 ;
        RECT 111.355 1.195 111.685 1.525 ;
        RECT 111.355 -0.165 111.685 0.165 ;
        RECT 111.36 -8.32 111.68 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.715 10.715 113.045 11.045 ;
        RECT 112.715 9.355 113.045 9.685 ;
        RECT 112.715 7.995 113.045 8.325 ;
        RECT 112.715 6.635 113.045 6.965 ;
        RECT 112.715 5.275 113.045 5.605 ;
        RECT 112.715 3.915 113.045 4.245 ;
        RECT 112.715 2.555 113.045 2.885 ;
        RECT 112.715 1.195 113.045 1.525 ;
        RECT 112.715 -0.165 113.045 0.165 ;
        RECT 112.72 -8.32 113.04 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.075 10.715 114.405 11.045 ;
        RECT 114.075 9.355 114.405 9.685 ;
        RECT 114.075 7.995 114.405 8.325 ;
        RECT 114.075 6.635 114.405 6.965 ;
        RECT 114.075 5.275 114.405 5.605 ;
        RECT 114.075 3.915 114.405 4.245 ;
        RECT 114.075 2.555 114.405 2.885 ;
        RECT 114.075 1.195 114.405 1.525 ;
        RECT 114.075 -0.165 114.405 0.165 ;
        RECT 114.08 -8.32 114.4 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.435 10.715 115.765 11.045 ;
        RECT 115.435 9.355 115.765 9.685 ;
        RECT 115.435 7.995 115.765 8.325 ;
        RECT 115.435 6.635 115.765 6.965 ;
        RECT 115.435 5.275 115.765 5.605 ;
        RECT 115.435 3.915 115.765 4.245 ;
        RECT 115.435 2.555 115.765 2.885 ;
        RECT 115.435 1.195 115.765 1.525 ;
        RECT 115.435 -0.165 115.765 0.165 ;
        RECT 115.44 -8.32 115.76 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.795 10.715 117.125 11.045 ;
        RECT 116.795 9.355 117.125 9.685 ;
        RECT 116.795 7.995 117.125 8.325 ;
        RECT 116.795 6.635 117.125 6.965 ;
        RECT 116.795 5.275 117.125 5.605 ;
        RECT 116.795 3.915 117.125 4.245 ;
        RECT 116.795 2.555 117.125 2.885 ;
        RECT 116.795 1.195 117.125 1.525 ;
        RECT 116.795 -0.165 117.125 0.165 ;
        RECT 116.8 -8.32 117.12 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.155 10.715 118.485 11.045 ;
        RECT 118.155 9.355 118.485 9.685 ;
        RECT 118.155 7.995 118.485 8.325 ;
        RECT 118.155 6.635 118.485 6.965 ;
        RECT 118.155 5.275 118.485 5.605 ;
        RECT 118.155 3.915 118.485 4.245 ;
        RECT 118.155 2.555 118.485 2.885 ;
        RECT 118.155 1.195 118.485 1.525 ;
        RECT 118.155 -0.165 118.485 0.165 ;
        RECT 118.16 -8.32 118.48 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 119.515 10.715 119.845 11.045 ;
        RECT 119.515 9.355 119.845 9.685 ;
        RECT 119.515 7.995 119.845 8.325 ;
        RECT 119.515 6.635 119.845 6.965 ;
        RECT 119.515 5.275 119.845 5.605 ;
        RECT 119.515 3.915 119.845 4.245 ;
        RECT 119.515 2.555 119.845 2.885 ;
        RECT 119.515 1.195 119.845 1.525 ;
        RECT 119.515 -0.165 119.845 0.165 ;
        RECT 119.52 -8.32 119.84 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.875 10.715 121.205 11.045 ;
        RECT 120.875 9.355 121.205 9.685 ;
        RECT 120.875 7.995 121.205 8.325 ;
        RECT 120.875 6.635 121.205 6.965 ;
        RECT 120.875 5.275 121.205 5.605 ;
        RECT 120.875 3.915 121.205 4.245 ;
        RECT 120.875 2.555 121.205 2.885 ;
        RECT 120.875 1.195 121.205 1.525 ;
        RECT 120.875 -0.165 121.205 0.165 ;
        RECT 120.88 -8.32 121.2 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.235 10.715 122.565 11.045 ;
        RECT 122.235 9.355 122.565 9.685 ;
        RECT 122.235 7.995 122.565 8.325 ;
        RECT 122.235 6.635 122.565 6.965 ;
        RECT 122.235 5.275 122.565 5.605 ;
        RECT 122.235 3.915 122.565 4.245 ;
        RECT 122.235 2.555 122.565 2.885 ;
        RECT 122.235 1.195 122.565 1.525 ;
        RECT 122.235 -0.165 122.565 0.165 ;
        RECT 122.24 -8.32 122.56 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.595 10.715 123.925 11.045 ;
        RECT 123.595 9.355 123.925 9.685 ;
        RECT 123.595 7.995 123.925 8.325 ;
        RECT 123.595 6.635 123.925 6.965 ;
        RECT 123.595 5.275 123.925 5.605 ;
        RECT 123.595 3.915 123.925 4.245 ;
        RECT 123.595 2.555 123.925 2.885 ;
        RECT 123.595 1.195 123.925 1.525 ;
        RECT 123.595 -0.165 123.925 0.165 ;
        RECT 123.6 -8.32 123.92 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.955 10.715 125.285 11.045 ;
        RECT 124.955 9.355 125.285 9.685 ;
        RECT 124.955 7.995 125.285 8.325 ;
        RECT 124.955 6.635 125.285 6.965 ;
        RECT 124.955 5.275 125.285 5.605 ;
        RECT 124.955 3.915 125.285 4.245 ;
        RECT 124.955 2.555 125.285 2.885 ;
        RECT 124.955 1.195 125.285 1.525 ;
        RECT 124.955 -0.165 125.285 0.165 ;
        RECT 124.96 -8.32 125.28 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.315 10.715 126.645 11.045 ;
        RECT 126.315 9.355 126.645 9.685 ;
        RECT 126.315 7.995 126.645 8.325 ;
        RECT 126.315 6.635 126.645 6.965 ;
        RECT 126.315 5.275 126.645 5.605 ;
        RECT 126.315 3.915 126.645 4.245 ;
        RECT 126.315 2.555 126.645 2.885 ;
        RECT 126.315 1.195 126.645 1.525 ;
        RECT 126.315 -0.165 126.645 0.165 ;
        RECT 126.32 -8.32 126.64 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.675 10.715 128.005 11.045 ;
        RECT 127.675 9.355 128.005 9.685 ;
        RECT 127.675 7.995 128.005 8.325 ;
        RECT 127.675 6.635 128.005 6.965 ;
        RECT 127.675 5.275 128.005 5.605 ;
        RECT 127.675 3.915 128.005 4.245 ;
        RECT 127.675 2.555 128.005 2.885 ;
        RECT 127.675 1.195 128.005 1.525 ;
        RECT 127.675 -0.165 128.005 0.165 ;
        RECT 127.68 -8.32 128 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.035 10.715 129.365 11.045 ;
        RECT 129.035 9.355 129.365 9.685 ;
        RECT 129.035 7.995 129.365 8.325 ;
        RECT 129.035 6.635 129.365 6.965 ;
        RECT 129.035 5.275 129.365 5.605 ;
        RECT 129.035 3.915 129.365 4.245 ;
        RECT 129.035 2.555 129.365 2.885 ;
        RECT 129.035 1.195 129.365 1.525 ;
        RECT 129.035 -0.165 129.365 0.165 ;
        RECT 129.04 -8.32 129.36 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.395 10.715 130.725 11.045 ;
        RECT 130.395 9.355 130.725 9.685 ;
        RECT 130.395 7.995 130.725 8.325 ;
        RECT 130.395 6.635 130.725 6.965 ;
        RECT 130.395 5.275 130.725 5.605 ;
        RECT 130.395 3.915 130.725 4.245 ;
        RECT 130.395 2.555 130.725 2.885 ;
        RECT 130.395 1.195 130.725 1.525 ;
        RECT 130.395 -0.165 130.725 0.165 ;
        RECT 130.4 -8.32 130.72 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.755 10.715 132.085 11.045 ;
        RECT 131.755 9.355 132.085 9.685 ;
        RECT 131.755 7.995 132.085 8.325 ;
        RECT 131.755 6.635 132.085 6.965 ;
        RECT 131.755 5.275 132.085 5.605 ;
        RECT 131.755 3.915 132.085 4.245 ;
        RECT 131.755 2.555 132.085 2.885 ;
        RECT 131.755 1.195 132.085 1.525 ;
        RECT 131.755 -0.165 132.085 0.165 ;
        RECT 131.76 -8.32 132.08 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.115 10.715 133.445 11.045 ;
        RECT 133.115 9.355 133.445 9.685 ;
        RECT 133.115 7.995 133.445 8.325 ;
        RECT 133.115 6.635 133.445 6.965 ;
        RECT 133.115 5.275 133.445 5.605 ;
        RECT 133.115 3.915 133.445 4.245 ;
        RECT 133.115 2.555 133.445 2.885 ;
        RECT 133.115 1.195 133.445 1.525 ;
        RECT 133.115 -0.165 133.445 0.165 ;
        RECT 133.12 -8.32 133.44 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.475 10.715 134.805 11.045 ;
        RECT 134.475 9.355 134.805 9.685 ;
        RECT 134.475 7.995 134.805 8.325 ;
        RECT 134.475 6.635 134.805 6.965 ;
        RECT 134.475 5.275 134.805 5.605 ;
        RECT 134.475 3.915 134.805 4.245 ;
        RECT 134.475 2.555 134.805 2.885 ;
        RECT 134.475 1.195 134.805 1.525 ;
        RECT 134.475 -0.165 134.805 0.165 ;
        RECT 134.48 -8.32 134.8 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.835 10.715 136.165 11.045 ;
        RECT 135.835 9.355 136.165 9.685 ;
        RECT 135.835 7.995 136.165 8.325 ;
        RECT 135.835 6.635 136.165 6.965 ;
        RECT 135.835 5.275 136.165 5.605 ;
        RECT 135.835 3.915 136.165 4.245 ;
        RECT 135.835 2.555 136.165 2.885 ;
        RECT 135.835 1.195 136.165 1.525 ;
        RECT 135.835 -0.165 136.165 0.165 ;
        RECT 135.84 -8.32 136.16 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.195 10.715 137.525 11.045 ;
        RECT 137.195 9.355 137.525 9.685 ;
        RECT 137.195 7.995 137.525 8.325 ;
        RECT 137.195 6.635 137.525 6.965 ;
        RECT 137.195 5.275 137.525 5.605 ;
        RECT 137.195 3.915 137.525 4.245 ;
        RECT 137.195 2.555 137.525 2.885 ;
        RECT 137.195 1.195 137.525 1.525 ;
        RECT 137.195 -0.165 137.525 0.165 ;
        RECT 137.2 -8.32 137.52 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 138.555 10.715 138.885 11.045 ;
        RECT 138.555 9.355 138.885 9.685 ;
        RECT 138.555 7.995 138.885 8.325 ;
        RECT 138.555 6.635 138.885 6.965 ;
        RECT 138.555 5.275 138.885 5.605 ;
        RECT 138.555 3.915 138.885 4.245 ;
        RECT 138.555 2.555 138.885 2.885 ;
        RECT 138.555 1.195 138.885 1.525 ;
        RECT 138.555 -0.165 138.885 0.165 ;
        RECT 138.56 -8.32 138.88 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.915 10.715 140.245 11.045 ;
        RECT 139.915 9.355 140.245 9.685 ;
        RECT 139.915 7.995 140.245 8.325 ;
        RECT 139.915 6.635 140.245 6.965 ;
        RECT 139.915 5.275 140.245 5.605 ;
        RECT 139.915 3.915 140.245 4.245 ;
        RECT 139.915 2.555 140.245 2.885 ;
        RECT 139.915 1.195 140.245 1.525 ;
        RECT 139.915 -0.165 140.245 0.165 ;
        RECT 139.92 -8.32 140.24 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.275 10.715 141.605 11.045 ;
        RECT 141.275 9.355 141.605 9.685 ;
        RECT 141.275 7.995 141.605 8.325 ;
        RECT 141.275 6.635 141.605 6.965 ;
        RECT 141.275 5.275 141.605 5.605 ;
        RECT 141.275 3.915 141.605 4.245 ;
        RECT 141.275 2.555 141.605 2.885 ;
        RECT 141.275 1.195 141.605 1.525 ;
        RECT 141.275 -0.165 141.605 0.165 ;
        RECT 141.28 -8.32 141.6 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.635 10.715 142.965 11.045 ;
        RECT 142.635 9.355 142.965 9.685 ;
        RECT 142.635 7.995 142.965 8.325 ;
        RECT 142.635 6.635 142.965 6.965 ;
        RECT 142.635 5.275 142.965 5.605 ;
        RECT 142.635 3.915 142.965 4.245 ;
        RECT 142.635 2.555 142.965 2.885 ;
        RECT 142.635 1.195 142.965 1.525 ;
        RECT 142.635 -0.165 142.965 0.165 ;
        RECT 142.64 -8.32 142.96 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.995 10.715 144.325 11.045 ;
        RECT 143.995 9.355 144.325 9.685 ;
        RECT 143.995 7.995 144.325 8.325 ;
        RECT 143.995 6.635 144.325 6.965 ;
        RECT 143.995 5.275 144.325 5.605 ;
        RECT 143.995 3.915 144.325 4.245 ;
        RECT 143.995 2.555 144.325 2.885 ;
        RECT 143.995 1.195 144.325 1.525 ;
        RECT 143.995 -0.165 144.325 0.165 ;
        RECT 144 -8.32 144.32 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.355 10.715 145.685 11.045 ;
        RECT 145.355 9.355 145.685 9.685 ;
        RECT 145.355 7.995 145.685 8.325 ;
        RECT 145.355 6.635 145.685 6.965 ;
        RECT 145.355 5.275 145.685 5.605 ;
        RECT 145.355 3.915 145.685 4.245 ;
        RECT 145.355 2.555 145.685 2.885 ;
        RECT 145.355 1.195 145.685 1.525 ;
        RECT 145.355 -0.165 145.685 0.165 ;
        RECT 145.36 -8.32 145.68 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.715 10.715 147.045 11.045 ;
        RECT 146.715 9.355 147.045 9.685 ;
        RECT 146.715 7.995 147.045 8.325 ;
        RECT 146.715 6.635 147.045 6.965 ;
        RECT 146.715 5.275 147.045 5.605 ;
        RECT 146.715 3.915 147.045 4.245 ;
        RECT 146.715 2.555 147.045 2.885 ;
        RECT 146.715 1.195 147.045 1.525 ;
        RECT 146.715 -0.165 147.045 0.165 ;
        RECT 146.72 -8.32 147.04 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.075 10.715 148.405 11.045 ;
        RECT 148.075 9.355 148.405 9.685 ;
        RECT 148.075 7.995 148.405 8.325 ;
        RECT 148.075 6.635 148.405 6.965 ;
        RECT 148.075 5.275 148.405 5.605 ;
        RECT 148.075 3.915 148.405 4.245 ;
        RECT 148.075 2.555 148.405 2.885 ;
        RECT 148.075 1.195 148.405 1.525 ;
        RECT 148.075 -0.165 148.405 0.165 ;
        RECT 148.08 -8.32 148.4 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.435 10.715 149.765 11.045 ;
        RECT 149.435 9.355 149.765 9.685 ;
        RECT 149.435 7.995 149.765 8.325 ;
        RECT 149.435 6.635 149.765 6.965 ;
        RECT 149.435 5.275 149.765 5.605 ;
        RECT 149.435 3.915 149.765 4.245 ;
        RECT 149.435 2.555 149.765 2.885 ;
        RECT 149.435 1.195 149.765 1.525 ;
        RECT 149.435 -0.165 149.765 0.165 ;
        RECT 149.44 -8.32 149.76 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.795 10.715 151.125 11.045 ;
        RECT 150.795 9.355 151.125 9.685 ;
        RECT 150.795 7.995 151.125 8.325 ;
        RECT 150.795 6.635 151.125 6.965 ;
        RECT 150.795 5.275 151.125 5.605 ;
        RECT 150.795 3.915 151.125 4.245 ;
        RECT 150.795 2.555 151.125 2.885 ;
        RECT 150.795 1.195 151.125 1.525 ;
        RECT 150.795 -0.165 151.125 0.165 ;
        RECT 150.8 -8.32 151.12 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.155 10.715 152.485 11.045 ;
        RECT 152.155 9.355 152.485 9.685 ;
        RECT 152.155 7.995 152.485 8.325 ;
        RECT 152.155 6.635 152.485 6.965 ;
        RECT 152.155 5.275 152.485 5.605 ;
        RECT 152.155 3.915 152.485 4.245 ;
        RECT 152.155 2.555 152.485 2.885 ;
        RECT 152.155 1.195 152.485 1.525 ;
        RECT 152.155 -0.165 152.485 0.165 ;
        RECT 152.16 -8.32 152.48 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.515 10.715 153.845 11.045 ;
        RECT 153.515 9.355 153.845 9.685 ;
        RECT 153.515 7.995 153.845 8.325 ;
        RECT 153.515 6.635 153.845 6.965 ;
        RECT 153.515 5.275 153.845 5.605 ;
        RECT 153.515 3.915 153.845 4.245 ;
        RECT 153.515 2.555 153.845 2.885 ;
        RECT 153.515 1.195 153.845 1.525 ;
        RECT 153.515 -0.165 153.845 0.165 ;
        RECT 153.52 -8.32 153.84 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.875 10.715 155.205 11.045 ;
        RECT 154.875 9.355 155.205 9.685 ;
        RECT 154.875 7.995 155.205 8.325 ;
        RECT 154.875 6.635 155.205 6.965 ;
        RECT 154.875 5.275 155.205 5.605 ;
        RECT 154.875 3.915 155.205 4.245 ;
        RECT 154.875 2.555 155.205 2.885 ;
        RECT 154.875 1.195 155.205 1.525 ;
        RECT 154.875 -0.165 155.205 0.165 ;
        RECT 154.88 -8.32 155.2 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.235 10.715 156.565 11.045 ;
        RECT 156.235 9.355 156.565 9.685 ;
        RECT 156.235 7.995 156.565 8.325 ;
        RECT 156.235 6.635 156.565 6.965 ;
        RECT 156.235 5.275 156.565 5.605 ;
        RECT 156.235 3.915 156.565 4.245 ;
        RECT 156.235 2.555 156.565 2.885 ;
        RECT 156.235 1.195 156.565 1.525 ;
        RECT 156.235 -0.165 156.565 0.165 ;
        RECT 156.24 -8.32 156.56 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 157.595 10.715 157.925 11.045 ;
        RECT 157.595 9.355 157.925 9.685 ;
        RECT 157.595 7.995 157.925 8.325 ;
        RECT 157.595 6.635 157.925 6.965 ;
        RECT 157.595 5.275 157.925 5.605 ;
        RECT 157.595 3.915 157.925 4.245 ;
        RECT 157.595 2.555 157.925 2.885 ;
        RECT 157.595 1.195 157.925 1.525 ;
        RECT 157.595 -0.165 157.925 0.165 ;
        RECT 157.6 -8.32 157.92 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.955 10.715 159.285 11.045 ;
        RECT 158.955 9.355 159.285 9.685 ;
        RECT 158.955 7.995 159.285 8.325 ;
        RECT 158.955 6.635 159.285 6.965 ;
        RECT 158.955 5.275 159.285 5.605 ;
        RECT 158.955 3.915 159.285 4.245 ;
        RECT 158.955 2.555 159.285 2.885 ;
        RECT 158.955 1.195 159.285 1.525 ;
        RECT 158.955 -0.165 159.285 0.165 ;
        RECT 158.96 -8.32 159.28 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.315 10.715 160.645 11.045 ;
        RECT 160.315 9.355 160.645 9.685 ;
        RECT 160.315 7.995 160.645 8.325 ;
        RECT 160.315 6.635 160.645 6.965 ;
        RECT 160.315 5.275 160.645 5.605 ;
        RECT 160.315 3.915 160.645 4.245 ;
        RECT 160.315 2.555 160.645 2.885 ;
        RECT 160.315 1.195 160.645 1.525 ;
        RECT 160.315 -0.165 160.645 0.165 ;
        RECT 160.32 -8.32 160.64 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.675 10.715 162.005 11.045 ;
        RECT 161.675 9.355 162.005 9.685 ;
        RECT 161.675 7.995 162.005 8.325 ;
        RECT 161.675 6.635 162.005 6.965 ;
        RECT 161.675 5.275 162.005 5.605 ;
        RECT 161.675 3.915 162.005 4.245 ;
        RECT 161.675 2.555 162.005 2.885 ;
        RECT 161.675 1.195 162.005 1.525 ;
        RECT 161.675 -0.165 162.005 0.165 ;
        RECT 161.68 -8.32 162 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.035 10.715 163.365 11.045 ;
        RECT 163.035 9.355 163.365 9.685 ;
        RECT 163.035 7.995 163.365 8.325 ;
        RECT 163.035 6.635 163.365 6.965 ;
        RECT 163.035 5.275 163.365 5.605 ;
        RECT 163.035 3.915 163.365 4.245 ;
        RECT 163.035 2.555 163.365 2.885 ;
        RECT 163.035 1.195 163.365 1.525 ;
        RECT 163.035 -0.165 163.365 0.165 ;
        RECT 163.04 -8.32 163.36 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 164.395 10.715 164.725 11.045 ;
        RECT 164.395 9.355 164.725 9.685 ;
        RECT 164.395 7.995 164.725 8.325 ;
        RECT 164.395 6.635 164.725 6.965 ;
        RECT 164.395 5.275 164.725 5.605 ;
        RECT 164.395 3.915 164.725 4.245 ;
        RECT 164.395 2.555 164.725 2.885 ;
        RECT 164.395 1.195 164.725 1.525 ;
        RECT 164.395 -0.165 164.725 0.165 ;
        RECT 164.4 -8.32 164.72 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.755 10.715 166.085 11.045 ;
        RECT 165.755 9.355 166.085 9.685 ;
        RECT 165.755 7.995 166.085 8.325 ;
        RECT 165.755 6.635 166.085 6.965 ;
        RECT 165.755 5.275 166.085 5.605 ;
        RECT 165.755 3.915 166.085 4.245 ;
        RECT 165.755 2.555 166.085 2.885 ;
        RECT 165.755 1.195 166.085 1.525 ;
        RECT 165.755 -0.165 166.085 0.165 ;
        RECT 165.76 -8.32 166.08 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.115 10.715 167.445 11.045 ;
        RECT 167.115 9.355 167.445 9.685 ;
        RECT 167.115 7.995 167.445 8.325 ;
        RECT 167.115 6.635 167.445 6.965 ;
        RECT 167.115 5.275 167.445 5.605 ;
        RECT 167.115 3.915 167.445 4.245 ;
        RECT 167.115 2.555 167.445 2.885 ;
        RECT 167.115 1.195 167.445 1.525 ;
        RECT 167.115 -0.165 167.445 0.165 ;
        RECT 167.12 -8.32 167.44 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 168.475 10.715 168.805 11.045 ;
        RECT 168.475 9.355 168.805 9.685 ;
        RECT 168.475 7.995 168.805 8.325 ;
        RECT 168.475 6.635 168.805 6.965 ;
        RECT 168.475 5.275 168.805 5.605 ;
        RECT 168.475 3.915 168.805 4.245 ;
        RECT 168.475 2.555 168.805 2.885 ;
        RECT 168.475 1.195 168.805 1.525 ;
        RECT 168.475 -0.165 168.805 0.165 ;
        RECT 168.48 -8.32 168.8 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.835 10.715 170.165 11.045 ;
        RECT 169.835 9.355 170.165 9.685 ;
        RECT 169.835 7.995 170.165 8.325 ;
        RECT 169.835 6.635 170.165 6.965 ;
        RECT 169.835 5.275 170.165 5.605 ;
        RECT 169.835 3.915 170.165 4.245 ;
        RECT 169.835 2.555 170.165 2.885 ;
        RECT 169.835 1.195 170.165 1.525 ;
        RECT 169.835 -0.165 170.165 0.165 ;
        RECT 169.84 -8.32 170.16 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.195 10.715 171.525 11.045 ;
        RECT 171.195 9.355 171.525 9.685 ;
        RECT 171.195 7.995 171.525 8.325 ;
        RECT 171.195 6.635 171.525 6.965 ;
        RECT 171.195 5.275 171.525 5.605 ;
        RECT 171.195 3.915 171.525 4.245 ;
        RECT 171.195 2.555 171.525 2.885 ;
        RECT 171.195 1.195 171.525 1.525 ;
        RECT 171.195 -0.165 171.525 0.165 ;
        RECT 171.2 -8.32 171.52 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.555 10.715 172.885 11.045 ;
        RECT 172.555 9.355 172.885 9.685 ;
        RECT 172.555 7.995 172.885 8.325 ;
        RECT 172.555 6.635 172.885 6.965 ;
        RECT 172.555 5.275 172.885 5.605 ;
        RECT 172.555 3.915 172.885 4.245 ;
        RECT 172.555 2.555 172.885 2.885 ;
        RECT 172.555 1.195 172.885 1.525 ;
        RECT 172.555 -0.165 172.885 0.165 ;
        RECT 172.56 -8.32 172.88 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.915 10.715 174.245 11.045 ;
        RECT 173.915 9.355 174.245 9.685 ;
        RECT 173.915 7.995 174.245 8.325 ;
        RECT 173.915 6.635 174.245 6.965 ;
        RECT 173.915 5.275 174.245 5.605 ;
        RECT 173.915 3.915 174.245 4.245 ;
        RECT 173.915 2.555 174.245 2.885 ;
        RECT 173.915 1.195 174.245 1.525 ;
        RECT 173.915 -0.165 174.245 0.165 ;
        RECT 173.92 -8.32 174.24 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.275 10.715 175.605 11.045 ;
        RECT 175.275 9.355 175.605 9.685 ;
        RECT 175.275 7.995 175.605 8.325 ;
        RECT 175.275 6.635 175.605 6.965 ;
        RECT 175.275 5.275 175.605 5.605 ;
        RECT 175.275 3.915 175.605 4.245 ;
        RECT 175.275 2.555 175.605 2.885 ;
        RECT 175.275 1.195 175.605 1.525 ;
        RECT 175.275 -0.165 175.605 0.165 ;
        RECT 175.28 -8.32 175.6 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 176.635 10.715 176.965 11.045 ;
        RECT 176.635 9.355 176.965 9.685 ;
        RECT 176.635 7.995 176.965 8.325 ;
        RECT 176.635 6.635 176.965 6.965 ;
        RECT 176.635 5.275 176.965 5.605 ;
        RECT 176.635 3.915 176.965 4.245 ;
        RECT 176.635 2.555 176.965 2.885 ;
        RECT 176.635 1.195 176.965 1.525 ;
        RECT 176.635 -0.165 176.965 0.165 ;
        RECT 176.64 -8.32 176.96 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.995 10.715 178.325 11.045 ;
        RECT 177.995 9.355 178.325 9.685 ;
        RECT 177.995 7.995 178.325 8.325 ;
        RECT 177.995 6.635 178.325 6.965 ;
        RECT 177.995 5.275 178.325 5.605 ;
        RECT 177.995 3.915 178.325 4.245 ;
        RECT 177.995 2.555 178.325 2.885 ;
        RECT 177.995 1.195 178.325 1.525 ;
        RECT 177.995 -0.165 178.325 0.165 ;
        RECT 178 -8.32 178.32 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 179.355 10.715 179.685 11.045 ;
        RECT 179.355 9.355 179.685 9.685 ;
        RECT 179.355 7.995 179.685 8.325 ;
        RECT 179.355 6.635 179.685 6.965 ;
        RECT 179.355 5.275 179.685 5.605 ;
        RECT 179.355 3.915 179.685 4.245 ;
        RECT 179.355 2.555 179.685 2.885 ;
        RECT 179.355 1.195 179.685 1.525 ;
        RECT 179.355 -0.165 179.685 0.165 ;
        RECT 179.36 -8.32 179.68 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.715 10.715 181.045 11.045 ;
        RECT 180.715 9.355 181.045 9.685 ;
        RECT 180.715 7.995 181.045 8.325 ;
        RECT 180.715 6.635 181.045 6.965 ;
        RECT 180.715 5.275 181.045 5.605 ;
        RECT 180.715 3.915 181.045 4.245 ;
        RECT 180.715 2.555 181.045 2.885 ;
        RECT 180.715 1.195 181.045 1.525 ;
        RECT 180.715 -0.165 181.045 0.165 ;
        RECT 180.72 -8.32 181.04 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.075 10.715 182.405 11.045 ;
        RECT 182.075 9.355 182.405 9.685 ;
        RECT 182.075 7.995 182.405 8.325 ;
        RECT 182.075 6.635 182.405 6.965 ;
        RECT 182.075 5.275 182.405 5.605 ;
        RECT 182.075 3.915 182.405 4.245 ;
        RECT 182.075 2.555 182.405 2.885 ;
        RECT 182.075 1.195 182.405 1.525 ;
        RECT 182.075 -0.165 182.405 0.165 ;
        RECT 182.08 -8.32 182.4 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 183.435 10.715 183.765 11.045 ;
        RECT 183.435 9.355 183.765 9.685 ;
        RECT 183.435 7.995 183.765 8.325 ;
        RECT 183.435 6.635 183.765 6.965 ;
        RECT 183.435 5.275 183.765 5.605 ;
        RECT 183.435 3.915 183.765 4.245 ;
        RECT 183.435 2.555 183.765 2.885 ;
        RECT 183.435 1.195 183.765 1.525 ;
        RECT 183.435 -0.165 183.765 0.165 ;
        RECT 183.44 -8.32 183.76 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.795 10.715 185.125 11.045 ;
        RECT 184.795 9.355 185.125 9.685 ;
        RECT 184.795 7.995 185.125 8.325 ;
        RECT 184.795 6.635 185.125 6.965 ;
        RECT 184.795 5.275 185.125 5.605 ;
        RECT 184.795 3.915 185.125 4.245 ;
        RECT 184.795 2.555 185.125 2.885 ;
        RECT 184.795 1.195 185.125 1.525 ;
        RECT 184.795 -0.165 185.125 0.165 ;
        RECT 184.8 -8.32 185.12 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.155 10.715 186.485 11.045 ;
        RECT 186.155 9.355 186.485 9.685 ;
        RECT 186.155 7.995 186.485 8.325 ;
        RECT 186.155 6.635 186.485 6.965 ;
        RECT 186.155 5.275 186.485 5.605 ;
        RECT 186.155 3.915 186.485 4.245 ;
        RECT 186.155 2.555 186.485 2.885 ;
        RECT 186.155 1.195 186.485 1.525 ;
        RECT 186.155 -0.165 186.485 0.165 ;
        RECT 186.16 -8.32 186.48 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 187.515 10.715 187.845 11.045 ;
        RECT 187.515 9.355 187.845 9.685 ;
        RECT 187.515 7.995 187.845 8.325 ;
        RECT 187.515 6.635 187.845 6.965 ;
        RECT 187.515 5.275 187.845 5.605 ;
        RECT 187.515 3.915 187.845 4.245 ;
        RECT 187.515 2.555 187.845 2.885 ;
        RECT 187.515 1.195 187.845 1.525 ;
        RECT 187.515 -0.165 187.845 0.165 ;
        RECT 187.52 -8.32 187.84 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.875 10.715 189.205 11.045 ;
        RECT 188.875 9.355 189.205 9.685 ;
        RECT 188.875 7.995 189.205 8.325 ;
        RECT 188.875 6.635 189.205 6.965 ;
        RECT 188.875 5.275 189.205 5.605 ;
        RECT 188.875 3.915 189.205 4.245 ;
        RECT 188.875 2.555 189.205 2.885 ;
        RECT 188.875 1.195 189.205 1.525 ;
        RECT 188.875 -0.165 189.205 0.165 ;
        RECT 188.88 -8.32 189.2 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.235 10.715 190.565 11.045 ;
        RECT 190.235 9.355 190.565 9.685 ;
        RECT 190.235 7.995 190.565 8.325 ;
        RECT 190.235 6.635 190.565 6.965 ;
        RECT 190.235 5.275 190.565 5.605 ;
        RECT 190.235 3.915 190.565 4.245 ;
        RECT 190.235 2.555 190.565 2.885 ;
        RECT 190.235 1.195 190.565 1.525 ;
        RECT 190.235 -0.165 190.565 0.165 ;
        RECT 190.24 -8.32 190.56 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 191.595 10.715 191.925 11.045 ;
        RECT 191.595 9.355 191.925 9.685 ;
        RECT 191.595 7.995 191.925 8.325 ;
        RECT 191.595 6.635 191.925 6.965 ;
        RECT 191.595 5.275 191.925 5.605 ;
        RECT 191.595 3.915 191.925 4.245 ;
        RECT 191.595 2.555 191.925 2.885 ;
        RECT 191.595 1.195 191.925 1.525 ;
        RECT 191.595 -0.165 191.925 0.165 ;
        RECT 191.6 -8.32 191.92 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.955 10.715 193.285 11.045 ;
        RECT 192.955 9.355 193.285 9.685 ;
        RECT 192.955 7.995 193.285 8.325 ;
        RECT 192.955 6.635 193.285 6.965 ;
        RECT 192.955 5.275 193.285 5.605 ;
        RECT 192.955 3.915 193.285 4.245 ;
        RECT 192.955 2.555 193.285 2.885 ;
        RECT 192.955 1.195 193.285 1.525 ;
        RECT 192.955 -0.165 193.285 0.165 ;
        RECT 192.96 -8.32 193.28 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.315 10.715 194.645 11.045 ;
        RECT 194.315 9.355 194.645 9.685 ;
        RECT 194.315 7.995 194.645 8.325 ;
        RECT 194.315 6.635 194.645 6.965 ;
        RECT 194.315 5.275 194.645 5.605 ;
        RECT 194.315 3.915 194.645 4.245 ;
        RECT 194.315 2.555 194.645 2.885 ;
        RECT 194.315 1.195 194.645 1.525 ;
        RECT 194.315 -0.165 194.645 0.165 ;
        RECT 194.32 -8.32 194.64 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 195.675 10.715 196.005 11.045 ;
        RECT 195.675 9.355 196.005 9.685 ;
        RECT 195.675 7.995 196.005 8.325 ;
        RECT 195.675 6.635 196.005 6.965 ;
        RECT 195.675 5.275 196.005 5.605 ;
        RECT 195.675 3.915 196.005 4.245 ;
        RECT 195.675 2.555 196.005 2.885 ;
        RECT 195.675 1.195 196.005 1.525 ;
        RECT 195.675 -0.165 196.005 0.165 ;
        RECT 195.68 -8.32 196 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.035 10.715 197.365 11.045 ;
        RECT 197.035 9.355 197.365 9.685 ;
        RECT 197.035 7.995 197.365 8.325 ;
        RECT 197.035 6.635 197.365 6.965 ;
        RECT 197.035 5.275 197.365 5.605 ;
        RECT 197.035 3.915 197.365 4.245 ;
        RECT 197.035 2.555 197.365 2.885 ;
        RECT 197.035 1.195 197.365 1.525 ;
        RECT 197.035 -0.165 197.365 0.165 ;
        RECT 197.04 -8.32 197.36 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.395 10.715 198.725 11.045 ;
        RECT 198.395 9.355 198.725 9.685 ;
        RECT 198.395 7.995 198.725 8.325 ;
        RECT 198.395 6.635 198.725 6.965 ;
        RECT 198.395 5.275 198.725 5.605 ;
        RECT 198.395 3.915 198.725 4.245 ;
        RECT 198.395 2.555 198.725 2.885 ;
        RECT 198.395 1.195 198.725 1.525 ;
        RECT 198.395 -0.165 198.725 0.165 ;
        RECT 198.4 -8.32 198.72 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.755 10.715 200.085 11.045 ;
        RECT 199.755 9.355 200.085 9.685 ;
        RECT 199.755 7.995 200.085 8.325 ;
        RECT 199.755 6.635 200.085 6.965 ;
        RECT 199.755 5.275 200.085 5.605 ;
        RECT 199.755 3.915 200.085 4.245 ;
        RECT 199.755 2.555 200.085 2.885 ;
        RECT 199.755 1.195 200.085 1.525 ;
        RECT 199.755 -0.165 200.085 0.165 ;
        RECT 199.76 -8.32 200.08 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.115 10.715 201.445 11.045 ;
        RECT 201.115 9.355 201.445 9.685 ;
        RECT 201.115 7.995 201.445 8.325 ;
        RECT 201.115 6.635 201.445 6.965 ;
        RECT 201.115 5.275 201.445 5.605 ;
        RECT 201.115 3.915 201.445 4.245 ;
        RECT 201.115 2.555 201.445 2.885 ;
        RECT 201.115 1.195 201.445 1.525 ;
        RECT 201.115 -0.165 201.445 0.165 ;
        RECT 201.12 -8.32 201.44 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 202.475 10.715 202.805 11.045 ;
        RECT 202.475 9.355 202.805 9.685 ;
        RECT 202.475 7.995 202.805 8.325 ;
        RECT 202.475 6.635 202.805 6.965 ;
        RECT 202.475 5.275 202.805 5.605 ;
        RECT 202.475 3.915 202.805 4.245 ;
        RECT 202.475 2.555 202.805 2.885 ;
        RECT 202.475 1.195 202.805 1.525 ;
        RECT 202.475 -0.165 202.805 0.165 ;
        RECT 202.48 -8.32 202.8 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.835 10.715 204.165 11.045 ;
        RECT 203.835 9.355 204.165 9.685 ;
        RECT 203.835 7.995 204.165 8.325 ;
        RECT 203.835 6.635 204.165 6.965 ;
        RECT 203.835 5.275 204.165 5.605 ;
        RECT 203.835 3.915 204.165 4.245 ;
        RECT 203.835 2.555 204.165 2.885 ;
        RECT 203.835 1.195 204.165 1.525 ;
        RECT 203.835 -0.165 204.165 0.165 ;
        RECT 203.84 -8.32 204.16 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.195 10.715 205.525 11.045 ;
        RECT 205.195 9.355 205.525 9.685 ;
        RECT 205.195 7.995 205.525 8.325 ;
        RECT 205.195 6.635 205.525 6.965 ;
        RECT 205.195 5.275 205.525 5.605 ;
        RECT 205.195 3.915 205.525 4.245 ;
        RECT 205.195 2.555 205.525 2.885 ;
        RECT 205.195 1.195 205.525 1.525 ;
        RECT 205.195 -0.165 205.525 0.165 ;
        RECT 205.2 -8.32 205.52 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 206.555 10.715 206.885 11.045 ;
        RECT 206.555 9.355 206.885 9.685 ;
        RECT 206.555 7.995 206.885 8.325 ;
        RECT 206.555 6.635 206.885 6.965 ;
        RECT 206.555 5.275 206.885 5.605 ;
        RECT 206.555 3.915 206.885 4.245 ;
        RECT 206.555 2.555 206.885 2.885 ;
        RECT 206.555 1.195 206.885 1.525 ;
        RECT 206.555 -0.165 206.885 0.165 ;
        RECT 206.56 -8.32 206.88 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.915 10.715 208.245 11.045 ;
        RECT 207.915 9.355 208.245 9.685 ;
        RECT 207.915 7.995 208.245 8.325 ;
        RECT 207.915 6.635 208.245 6.965 ;
        RECT 207.915 5.275 208.245 5.605 ;
        RECT 207.915 3.915 208.245 4.245 ;
        RECT 207.915 2.555 208.245 2.885 ;
        RECT 207.915 1.195 208.245 1.525 ;
        RECT 207.915 -0.165 208.245 0.165 ;
        RECT 207.92 -8.32 208.24 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.275 10.715 209.605 11.045 ;
        RECT 209.275 9.355 209.605 9.685 ;
        RECT 209.275 7.995 209.605 8.325 ;
        RECT 209.275 6.635 209.605 6.965 ;
        RECT 209.275 5.275 209.605 5.605 ;
        RECT 209.275 3.915 209.605 4.245 ;
        RECT 209.275 2.555 209.605 2.885 ;
        RECT 209.275 1.195 209.605 1.525 ;
        RECT 209.275 -0.165 209.605 0.165 ;
        RECT 209.28 -8.32 209.6 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 210.635 10.715 210.965 11.045 ;
        RECT 210.635 9.355 210.965 9.685 ;
        RECT 210.635 7.995 210.965 8.325 ;
        RECT 210.635 6.635 210.965 6.965 ;
        RECT 210.635 5.275 210.965 5.605 ;
        RECT 210.635 3.915 210.965 4.245 ;
        RECT 210.635 2.555 210.965 2.885 ;
        RECT 210.635 1.195 210.965 1.525 ;
        RECT 210.635 -0.165 210.965 0.165 ;
        RECT 210.64 -8.32 210.96 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 211.995 10.715 212.325 11.045 ;
        RECT 211.995 9.355 212.325 9.685 ;
        RECT 211.995 7.995 212.325 8.325 ;
        RECT 211.995 6.635 212.325 6.965 ;
        RECT 211.995 5.275 212.325 5.605 ;
        RECT 211.995 3.915 212.325 4.245 ;
        RECT 211.995 2.555 212.325 2.885 ;
        RECT 211.995 1.195 212.325 1.525 ;
        RECT 211.995 -0.165 212.325 0.165 ;
        RECT 212 -8.32 212.32 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 213.355 10.715 213.685 11.045 ;
        RECT 213.355 9.355 213.685 9.685 ;
        RECT 213.355 7.995 213.685 8.325 ;
        RECT 213.355 6.635 213.685 6.965 ;
        RECT 213.355 5.275 213.685 5.605 ;
        RECT 213.355 3.915 213.685 4.245 ;
        RECT 213.355 2.555 213.685 2.885 ;
        RECT 213.355 1.195 213.685 1.525 ;
        RECT 213.355 -0.165 213.685 0.165 ;
        RECT 213.36 -8.32 213.68 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.715 10.715 215.045 11.045 ;
        RECT 214.715 9.355 215.045 9.685 ;
        RECT 214.715 7.995 215.045 8.325 ;
        RECT 214.715 6.635 215.045 6.965 ;
        RECT 214.715 5.275 215.045 5.605 ;
        RECT 214.715 3.915 215.045 4.245 ;
        RECT 214.715 2.555 215.045 2.885 ;
        RECT 214.715 1.195 215.045 1.525 ;
        RECT 214.715 -0.165 215.045 0.165 ;
        RECT 214.72 -8.32 215.04 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.075 10.715 216.405 11.045 ;
        RECT 216.075 9.355 216.405 9.685 ;
        RECT 216.075 7.995 216.405 8.325 ;
        RECT 216.075 6.635 216.405 6.965 ;
        RECT 216.075 5.275 216.405 5.605 ;
        RECT 216.075 3.915 216.405 4.245 ;
        RECT 216.075 2.555 216.405 2.885 ;
        RECT 216.075 1.195 216.405 1.525 ;
        RECT 216.075 -0.165 216.405 0.165 ;
        RECT 216.08 -8.32 216.4 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 217.435 10.715 217.765 11.045 ;
        RECT 217.435 9.355 217.765 9.685 ;
        RECT 217.435 7.995 217.765 8.325 ;
        RECT 217.435 6.635 217.765 6.965 ;
        RECT 217.435 5.275 217.765 5.605 ;
        RECT 217.435 3.915 217.765 4.245 ;
        RECT 217.435 2.555 217.765 2.885 ;
        RECT 217.435 1.195 217.765 1.525 ;
        RECT 217.435 -0.165 217.765 0.165 ;
        RECT 217.44 -8.32 217.76 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.795 10.715 219.125 11.045 ;
        RECT 218.795 9.355 219.125 9.685 ;
        RECT 218.795 7.995 219.125 8.325 ;
        RECT 218.795 6.635 219.125 6.965 ;
        RECT 218.795 5.275 219.125 5.605 ;
        RECT 218.795 3.915 219.125 4.245 ;
        RECT 218.795 2.555 219.125 2.885 ;
        RECT 218.795 1.195 219.125 1.525 ;
        RECT 218.795 -0.165 219.125 0.165 ;
        RECT 218.8 -8.32 219.12 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.155 10.715 220.485 11.045 ;
        RECT 220.155 9.355 220.485 9.685 ;
        RECT 220.155 7.995 220.485 8.325 ;
        RECT 220.155 6.635 220.485 6.965 ;
        RECT 220.155 5.275 220.485 5.605 ;
        RECT 220.155 3.915 220.485 4.245 ;
        RECT 220.155 2.555 220.485 2.885 ;
        RECT 220.155 1.195 220.485 1.525 ;
        RECT 220.155 -0.165 220.485 0.165 ;
        RECT 220.16 -8.32 220.48 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 221.515 10.715 221.845 11.045 ;
        RECT 221.515 9.355 221.845 9.685 ;
        RECT 221.515 7.995 221.845 8.325 ;
        RECT 221.515 6.635 221.845 6.965 ;
        RECT 221.515 5.275 221.845 5.605 ;
        RECT 221.515 3.915 221.845 4.245 ;
        RECT 221.515 2.555 221.845 2.885 ;
        RECT 221.515 1.195 221.845 1.525 ;
        RECT 221.515 -0.165 221.845 0.165 ;
        RECT 221.52 -8.32 221.84 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.875 10.715 223.205 11.045 ;
        RECT 222.875 9.355 223.205 9.685 ;
        RECT 222.875 7.995 223.205 8.325 ;
        RECT 222.875 6.635 223.205 6.965 ;
        RECT 222.875 5.275 223.205 5.605 ;
        RECT 222.875 3.915 223.205 4.245 ;
        RECT 222.875 2.555 223.205 2.885 ;
        RECT 222.875 1.195 223.205 1.525 ;
        RECT 222.875 -0.165 223.205 0.165 ;
        RECT 222.88 -8.32 223.2 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 224.235 10.715 224.565 11.045 ;
        RECT 224.235 9.355 224.565 9.685 ;
        RECT 224.235 7.995 224.565 8.325 ;
        RECT 224.235 6.635 224.565 6.965 ;
        RECT 224.235 5.275 224.565 5.605 ;
        RECT 224.235 3.915 224.565 4.245 ;
        RECT 224.235 2.555 224.565 2.885 ;
        RECT 224.235 1.195 224.565 1.525 ;
        RECT 224.235 -0.165 224.565 0.165 ;
        RECT 224.24 -8.32 224.56 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 225.595 9.355 225.925 9.685 ;
        RECT 225.595 7.995 225.925 8.325 ;
        RECT 225.595 6.635 225.925 6.965 ;
        RECT 225.595 5.275 225.925 5.605 ;
        RECT 225.595 3.915 225.925 4.245 ;
        RECT 225.595 2.555 225.925 2.885 ;
        RECT 225.595 1.195 225.925 1.525 ;
        RECT 225.595 -0.165 225.925 0.165 ;
        RECT 225.6 -8.32 225.92 15.8 ;
        RECT 225.595 10.715 225.925 11.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -2.885 14.795 -2.555 15.125 ;
        RECT -2.885 13.435 -2.555 13.765 ;
        RECT -2.885 12.075 -2.555 12.405 ;
        RECT -2.885 10.715 -2.555 11.045 ;
        RECT -2.885 9.355 -2.555 9.685 ;
        RECT -2.885 7.995 -2.555 8.325 ;
        RECT -2.885 6.635 -2.555 6.965 ;
        RECT -2.885 5.275 -2.555 5.605 ;
        RECT -2.885 3.915 -2.555 4.245 ;
        RECT -2.885 2.555 -2.555 2.885 ;
        RECT -2.885 1.195 -2.555 1.525 ;
        RECT -2.885 -0.165 -2.555 0.165 ;
        RECT -2.88 -8.32 -2.56 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.525 14.795 -1.195 15.125 ;
        RECT -1.525 13.435 -1.195 13.765 ;
        RECT -1.525 12.075 -1.195 12.405 ;
        RECT -1.525 10.715 -1.195 11.045 ;
        RECT -1.525 9.355 -1.195 9.685 ;
        RECT -1.525 7.995 -1.195 8.325 ;
        RECT -1.525 6.635 -1.195 6.965 ;
        RECT -1.525 5.275 -1.195 5.605 ;
        RECT -1.525 3.915 -1.195 4.245 ;
        RECT -1.525 2.555 -1.195 2.885 ;
        RECT -1.525 1.195 -1.195 1.525 ;
        RECT -1.525 -0.165 -1.195 0.165 ;
        RECT -1.52 -8.32 -1.2 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.165 13.435 0.165 13.765 ;
        RECT -0.165 12.075 0.165 12.405 ;
        RECT -0.165 10.715 0.165 11.045 ;
        RECT -0.165 9.355 0.165 9.685 ;
        RECT -0.165 7.995 0.165 8.325 ;
        RECT -0.165 6.635 0.165 6.965 ;
        RECT -0.165 5.275 0.165 5.605 ;
        RECT -0.165 3.915 0.165 4.245 ;
        RECT -0.165 2.555 0.165 2.885 ;
        RECT -0.165 1.195 0.165 1.525 ;
        RECT -0.165 -0.165 0.165 0.165 ;
        RECT -0.16 -8.32 0.16 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.195 13.435 1.525 13.765 ;
        RECT 1.195 10.715 1.525 11.045 ;
        RECT 1.195 9.355 1.525 9.685 ;
        RECT 1.195 7.995 1.525 8.325 ;
        RECT 1.195 6.635 1.525 6.965 ;
        RECT 1.195 5.275 1.525 5.605 ;
        RECT 1.195 3.915 1.525 4.245 ;
        RECT 1.195 2.555 1.525 2.885 ;
        RECT 1.195 1.195 1.525 1.525 ;
        RECT 1.195 -0.165 1.525 0.165 ;
        RECT 1.2 -8.32 1.52 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 13.435 2.885 13.765 ;
        RECT 2.555 10.715 2.885 11.045 ;
        RECT 2.555 9.355 2.885 9.685 ;
        RECT 2.555 7.995 2.885 8.325 ;
        RECT 2.555 6.635 2.885 6.965 ;
        RECT 2.555 5.275 2.885 5.605 ;
        RECT 2.555 3.915 2.885 4.245 ;
        RECT 2.555 2.555 2.885 2.885 ;
        RECT 2.555 1.195 2.885 1.525 ;
        RECT 2.555 -0.165 2.885 0.165 ;
        RECT 2.56 -8.32 2.88 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.915 10.715 4.245 11.045 ;
        RECT 3.915 9.355 4.245 9.685 ;
        RECT 3.915 7.995 4.245 8.325 ;
        RECT 3.915 6.635 4.245 6.965 ;
        RECT 3.915 5.275 4.245 5.605 ;
        RECT 3.915 3.915 4.245 4.245 ;
        RECT 3.915 2.555 4.245 2.885 ;
        RECT 3.915 1.195 4.245 1.525 ;
        RECT 3.915 -0.165 4.245 0.165 ;
        RECT 3.92 -8.32 4.24 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.275 10.715 5.605 11.045 ;
        RECT 5.275 9.355 5.605 9.685 ;
        RECT 5.275 7.995 5.605 8.325 ;
        RECT 5.275 6.635 5.605 6.965 ;
        RECT 5.275 5.275 5.605 5.605 ;
        RECT 5.275 3.915 5.605 4.245 ;
        RECT 5.275 2.555 5.605 2.885 ;
        RECT 5.275 1.195 5.605 1.525 ;
        RECT 5.275 -0.165 5.605 0.165 ;
        RECT 5.28 -8.32 5.6 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 10.715 6.965 11.045 ;
        RECT 6.635 9.355 6.965 9.685 ;
        RECT 6.635 7.995 6.965 8.325 ;
        RECT 6.635 6.635 6.965 6.965 ;
        RECT 6.635 5.275 6.965 5.605 ;
        RECT 6.635 3.915 6.965 4.245 ;
        RECT 6.635 2.555 6.965 2.885 ;
        RECT 6.635 1.195 6.965 1.525 ;
        RECT 6.635 -0.165 6.965 0.165 ;
        RECT 6.64 -8.32 6.96 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.995 10.715 8.325 11.045 ;
        RECT 7.995 9.355 8.325 9.685 ;
        RECT 7.995 7.995 8.325 8.325 ;
        RECT 7.995 6.635 8.325 6.965 ;
        RECT 7.995 5.275 8.325 5.605 ;
        RECT 7.995 3.915 8.325 4.245 ;
        RECT 7.995 2.555 8.325 2.885 ;
        RECT 7.995 1.195 8.325 1.525 ;
        RECT 7.995 -0.165 8.325 0.165 ;
        RECT 8 -8.32 8.32 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 10.715 9.685 11.045 ;
        RECT 9.355 9.355 9.685 9.685 ;
        RECT 9.355 7.995 9.685 8.325 ;
        RECT 9.355 6.635 9.685 6.965 ;
        RECT 9.355 5.275 9.685 5.605 ;
        RECT 9.355 3.915 9.685 4.245 ;
        RECT 9.355 2.555 9.685 2.885 ;
        RECT 9.355 1.195 9.685 1.525 ;
        RECT 9.355 -0.165 9.685 0.165 ;
        RECT 9.36 -8.32 9.68 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.715 10.715 11.045 11.045 ;
        RECT 10.715 9.355 11.045 9.685 ;
        RECT 10.715 7.995 11.045 8.325 ;
        RECT 10.715 6.635 11.045 6.965 ;
        RECT 10.715 5.275 11.045 5.605 ;
        RECT 10.715 3.915 11.045 4.245 ;
        RECT 10.715 2.555 11.045 2.885 ;
        RECT 10.715 1.195 11.045 1.525 ;
        RECT 10.715 -0.165 11.045 0.165 ;
        RECT 10.72 -8.32 11.04 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.075 10.715 12.405 11.045 ;
        RECT 12.075 9.355 12.405 9.685 ;
        RECT 12.075 7.995 12.405 8.325 ;
        RECT 12.075 6.635 12.405 6.965 ;
        RECT 12.075 5.275 12.405 5.605 ;
        RECT 12.075 3.915 12.405 4.245 ;
        RECT 12.075 2.555 12.405 2.885 ;
        RECT 12.075 1.195 12.405 1.525 ;
        RECT 12.075 -0.165 12.405 0.165 ;
        RECT 12.08 -8.32 12.4 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.435 10.715 13.765 11.045 ;
        RECT 13.435 9.355 13.765 9.685 ;
        RECT 13.435 7.995 13.765 8.325 ;
        RECT 13.435 6.635 13.765 6.965 ;
        RECT 13.435 5.275 13.765 5.605 ;
        RECT 13.435 3.915 13.765 4.245 ;
        RECT 13.435 2.555 13.765 2.885 ;
        RECT 13.435 1.195 13.765 1.525 ;
        RECT 13.435 -0.165 13.765 0.165 ;
        RECT 13.44 -8.32 13.76 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.795 10.715 15.125 11.045 ;
        RECT 14.795 9.355 15.125 9.685 ;
        RECT 14.795 7.995 15.125 8.325 ;
        RECT 14.795 6.635 15.125 6.965 ;
        RECT 14.795 5.275 15.125 5.605 ;
        RECT 14.795 3.915 15.125 4.245 ;
        RECT 14.795 2.555 15.125 2.885 ;
        RECT 14.795 1.195 15.125 1.525 ;
        RECT 14.795 -0.165 15.125 0.165 ;
        RECT 14.8 -8.32 15.12 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.155 10.715 16.485 11.045 ;
        RECT 16.155 9.355 16.485 9.685 ;
        RECT 16.155 7.995 16.485 8.325 ;
        RECT 16.155 6.635 16.485 6.965 ;
        RECT 16.155 5.275 16.485 5.605 ;
        RECT 16.155 3.915 16.485 4.245 ;
        RECT 16.155 2.555 16.485 2.885 ;
        RECT 16.155 1.195 16.485 1.525 ;
        RECT 16.155 -0.165 16.485 0.165 ;
        RECT 16.16 -8.32 16.48 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.515 10.715 17.845 11.045 ;
        RECT 17.515 9.355 17.845 9.685 ;
        RECT 17.515 7.995 17.845 8.325 ;
        RECT 17.515 6.635 17.845 6.965 ;
        RECT 17.515 5.275 17.845 5.605 ;
        RECT 17.515 3.915 17.845 4.245 ;
        RECT 17.515 2.555 17.845 2.885 ;
        RECT 17.515 1.195 17.845 1.525 ;
        RECT 17.515 -0.165 17.845 0.165 ;
        RECT 17.52 -8.32 17.84 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.875 10.715 19.205 11.045 ;
        RECT 18.875 9.355 19.205 9.685 ;
        RECT 18.875 7.995 19.205 8.325 ;
        RECT 18.875 6.635 19.205 6.965 ;
        RECT 18.875 5.275 19.205 5.605 ;
        RECT 18.875 3.915 19.205 4.245 ;
        RECT 18.875 2.555 19.205 2.885 ;
        RECT 18.875 1.195 19.205 1.525 ;
        RECT 18.875 -0.165 19.205 0.165 ;
        RECT 18.88 -8.32 19.2 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.235 10.715 20.565 11.045 ;
        RECT 20.235 9.355 20.565 9.685 ;
        RECT 20.235 7.995 20.565 8.325 ;
        RECT 20.235 6.635 20.565 6.965 ;
        RECT 20.235 5.275 20.565 5.605 ;
        RECT 20.235 3.915 20.565 4.245 ;
        RECT 20.235 2.555 20.565 2.885 ;
        RECT 20.235 1.195 20.565 1.525 ;
        RECT 20.235 -0.165 20.565 0.165 ;
        RECT 20.24 -8.32 20.56 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.595 10.715 21.925 11.045 ;
        RECT 21.595 9.355 21.925 9.685 ;
        RECT 21.595 7.995 21.925 8.325 ;
        RECT 21.595 6.635 21.925 6.965 ;
        RECT 21.595 5.275 21.925 5.605 ;
        RECT 21.595 3.915 21.925 4.245 ;
        RECT 21.595 2.555 21.925 2.885 ;
        RECT 21.595 1.195 21.925 1.525 ;
        RECT 21.595 -0.165 21.925 0.165 ;
        RECT 21.6 -8.32 21.92 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.955 10.715 23.285 11.045 ;
        RECT 22.955 9.355 23.285 9.685 ;
        RECT 22.955 7.995 23.285 8.325 ;
        RECT 22.955 6.635 23.285 6.965 ;
        RECT 22.955 5.275 23.285 5.605 ;
        RECT 22.955 3.915 23.285 4.245 ;
        RECT 22.955 2.555 23.285 2.885 ;
        RECT 22.955 1.195 23.285 1.525 ;
        RECT 22.955 -0.165 23.285 0.165 ;
        RECT 22.96 -8.32 23.28 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.315 10.715 24.645 11.045 ;
        RECT 24.315 9.355 24.645 9.685 ;
        RECT 24.315 7.995 24.645 8.325 ;
        RECT 24.315 6.635 24.645 6.965 ;
        RECT 24.315 5.275 24.645 5.605 ;
        RECT 24.315 3.915 24.645 4.245 ;
        RECT 24.315 2.555 24.645 2.885 ;
        RECT 24.315 1.195 24.645 1.525 ;
        RECT 24.315 -0.165 24.645 0.165 ;
        RECT 24.32 -8.32 24.64 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.675 10.715 26.005 11.045 ;
        RECT 25.675 9.355 26.005 9.685 ;
        RECT 25.675 7.995 26.005 8.325 ;
        RECT 25.675 6.635 26.005 6.965 ;
        RECT 25.675 5.275 26.005 5.605 ;
        RECT 25.675 3.915 26.005 4.245 ;
        RECT 25.675 2.555 26.005 2.885 ;
        RECT 25.675 1.195 26.005 1.525 ;
        RECT 25.675 -0.165 26.005 0.165 ;
        RECT 25.68 -8.32 26 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.035 10.715 27.365 11.045 ;
        RECT 27.035 9.355 27.365 9.685 ;
        RECT 27.035 7.995 27.365 8.325 ;
        RECT 27.035 6.635 27.365 6.965 ;
        RECT 27.035 5.275 27.365 5.605 ;
        RECT 27.035 3.915 27.365 4.245 ;
        RECT 27.035 2.555 27.365 2.885 ;
        RECT 27.035 1.195 27.365 1.525 ;
        RECT 27.035 -0.165 27.365 0.165 ;
        RECT 27.04 -8.32 27.36 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.395 10.715 28.725 11.045 ;
        RECT 28.395 9.355 28.725 9.685 ;
        RECT 28.395 7.995 28.725 8.325 ;
        RECT 28.395 6.635 28.725 6.965 ;
        RECT 28.395 5.275 28.725 5.605 ;
        RECT 28.395 3.915 28.725 4.245 ;
        RECT 28.395 2.555 28.725 2.885 ;
        RECT 28.395 1.195 28.725 1.525 ;
        RECT 28.395 -0.165 28.725 0.165 ;
        RECT 28.4 -8.32 28.72 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.755 10.715 30.085 11.045 ;
        RECT 29.755 9.355 30.085 9.685 ;
        RECT 29.755 7.995 30.085 8.325 ;
        RECT 29.755 6.635 30.085 6.965 ;
        RECT 29.755 5.275 30.085 5.605 ;
        RECT 29.755 3.915 30.085 4.245 ;
        RECT 29.755 2.555 30.085 2.885 ;
        RECT 29.755 1.195 30.085 1.525 ;
        RECT 29.755 -0.165 30.085 0.165 ;
        RECT 29.76 -8.32 30.08 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.115 10.715 31.445 11.045 ;
        RECT 31.115 9.355 31.445 9.685 ;
        RECT 31.115 7.995 31.445 8.325 ;
        RECT 31.115 6.635 31.445 6.965 ;
        RECT 31.115 5.275 31.445 5.605 ;
        RECT 31.115 3.915 31.445 4.245 ;
        RECT 31.115 2.555 31.445 2.885 ;
        RECT 31.115 1.195 31.445 1.525 ;
        RECT 31.115 -0.165 31.445 0.165 ;
        RECT 31.12 -8.32 31.44 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.475 10.715 32.805 11.045 ;
        RECT 32.475 9.355 32.805 9.685 ;
        RECT 32.475 7.995 32.805 8.325 ;
        RECT 32.475 6.635 32.805 6.965 ;
        RECT 32.475 5.275 32.805 5.605 ;
        RECT 32.475 3.915 32.805 4.245 ;
        RECT 32.475 2.555 32.805 2.885 ;
        RECT 32.475 1.195 32.805 1.525 ;
        RECT 32.475 -0.165 32.805 0.165 ;
        RECT 32.48 -8.32 32.8 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.835 10.715 34.165 11.045 ;
        RECT 33.835 9.355 34.165 9.685 ;
        RECT 33.835 7.995 34.165 8.325 ;
        RECT 33.835 6.635 34.165 6.965 ;
        RECT 33.835 5.275 34.165 5.605 ;
        RECT 33.835 3.915 34.165 4.245 ;
        RECT 33.835 2.555 34.165 2.885 ;
        RECT 33.835 1.195 34.165 1.525 ;
        RECT 33.835 -0.165 34.165 0.165 ;
        RECT 33.84 -8.32 34.16 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.195 10.715 35.525 11.045 ;
        RECT 35.195 9.355 35.525 9.685 ;
        RECT 35.195 7.995 35.525 8.325 ;
        RECT 35.195 6.635 35.525 6.965 ;
        RECT 35.195 5.275 35.525 5.605 ;
        RECT 35.195 3.915 35.525 4.245 ;
        RECT 35.195 2.555 35.525 2.885 ;
        RECT 35.195 1.195 35.525 1.525 ;
        RECT 35.195 -0.165 35.525 0.165 ;
        RECT 35.2 -8.32 35.52 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.555 10.715 36.885 11.045 ;
        RECT 36.555 9.355 36.885 9.685 ;
        RECT 36.555 7.995 36.885 8.325 ;
        RECT 36.555 6.635 36.885 6.965 ;
        RECT 36.555 5.275 36.885 5.605 ;
        RECT 36.555 3.915 36.885 4.245 ;
        RECT 36.555 2.555 36.885 2.885 ;
        RECT 36.555 1.195 36.885 1.525 ;
        RECT 36.555 -0.165 36.885 0.165 ;
        RECT 36.56 -8.32 36.88 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.915 10.715 38.245 11.045 ;
        RECT 37.915 9.355 38.245 9.685 ;
        RECT 37.915 7.995 38.245 8.325 ;
        RECT 37.915 6.635 38.245 6.965 ;
        RECT 37.915 5.275 38.245 5.605 ;
        RECT 37.915 3.915 38.245 4.245 ;
        RECT 37.915 2.555 38.245 2.885 ;
        RECT 37.915 1.195 38.245 1.525 ;
        RECT 37.915 -0.165 38.245 0.165 ;
        RECT 37.92 -8.32 38.24 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.275 10.715 39.605 11.045 ;
        RECT 39.275 9.355 39.605 9.685 ;
        RECT 39.275 7.995 39.605 8.325 ;
        RECT 39.275 6.635 39.605 6.965 ;
        RECT 39.275 5.275 39.605 5.605 ;
        RECT 39.275 3.915 39.605 4.245 ;
        RECT 39.275 2.555 39.605 2.885 ;
        RECT 39.275 1.195 39.605 1.525 ;
        RECT 39.275 -0.165 39.605 0.165 ;
        RECT 39.28 -8.32 39.6 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.635 10.715 40.965 11.045 ;
        RECT 40.635 9.355 40.965 9.685 ;
        RECT 40.635 7.995 40.965 8.325 ;
        RECT 40.635 6.635 40.965 6.965 ;
        RECT 40.635 5.275 40.965 5.605 ;
        RECT 40.635 3.915 40.965 4.245 ;
        RECT 40.635 2.555 40.965 2.885 ;
        RECT 40.635 1.195 40.965 1.525 ;
        RECT 40.635 -0.165 40.965 0.165 ;
        RECT 40.64 -8.32 40.96 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.995 10.715 42.325 11.045 ;
        RECT 41.995 9.355 42.325 9.685 ;
        RECT 41.995 7.995 42.325 8.325 ;
        RECT 41.995 6.635 42.325 6.965 ;
        RECT 41.995 5.275 42.325 5.605 ;
        RECT 41.995 3.915 42.325 4.245 ;
        RECT 41.995 2.555 42.325 2.885 ;
        RECT 41.995 1.195 42.325 1.525 ;
        RECT 41.995 -0.165 42.325 0.165 ;
        RECT 42 -8.32 42.32 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.355 10.715 43.685 11.045 ;
        RECT 43.355 9.355 43.685 9.685 ;
        RECT 43.355 7.995 43.685 8.325 ;
        RECT 43.355 6.635 43.685 6.965 ;
        RECT 43.355 5.275 43.685 5.605 ;
        RECT 43.355 3.915 43.685 4.245 ;
        RECT 43.355 2.555 43.685 2.885 ;
        RECT 43.355 1.195 43.685 1.525 ;
        RECT 43.355 -0.165 43.685 0.165 ;
        RECT 43.36 -8.32 43.68 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.715 10.715 45.045 11.045 ;
        RECT 44.715 9.355 45.045 9.685 ;
        RECT 44.715 7.995 45.045 8.325 ;
        RECT 44.715 6.635 45.045 6.965 ;
        RECT 44.715 5.275 45.045 5.605 ;
        RECT 44.715 3.915 45.045 4.245 ;
        RECT 44.715 2.555 45.045 2.885 ;
        RECT 44.715 1.195 45.045 1.525 ;
        RECT 44.715 -0.165 45.045 0.165 ;
        RECT 44.72 -8.32 45.04 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.075 10.715 46.405 11.045 ;
        RECT 46.075 9.355 46.405 9.685 ;
        RECT 46.075 7.995 46.405 8.325 ;
        RECT 46.075 6.635 46.405 6.965 ;
        RECT 46.075 5.275 46.405 5.605 ;
        RECT 46.075 3.915 46.405 4.245 ;
        RECT 46.075 2.555 46.405 2.885 ;
        RECT 46.075 1.195 46.405 1.525 ;
        RECT 46.075 -0.165 46.405 0.165 ;
        RECT 46.08 -8.32 46.4 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.435 10.715 47.765 11.045 ;
        RECT 47.435 9.355 47.765 9.685 ;
        RECT 47.435 7.995 47.765 8.325 ;
        RECT 47.435 6.635 47.765 6.965 ;
        RECT 47.435 5.275 47.765 5.605 ;
        RECT 47.435 3.915 47.765 4.245 ;
        RECT 47.435 2.555 47.765 2.885 ;
        RECT 47.435 1.195 47.765 1.525 ;
        RECT 47.435 -0.165 47.765 0.165 ;
        RECT 47.44 -8.32 47.76 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.795 10.715 49.125 11.045 ;
        RECT 48.795 9.355 49.125 9.685 ;
        RECT 48.795 7.995 49.125 8.325 ;
        RECT 48.795 6.635 49.125 6.965 ;
        RECT 48.795 5.275 49.125 5.605 ;
        RECT 48.795 3.915 49.125 4.245 ;
        RECT 48.795 2.555 49.125 2.885 ;
        RECT 48.795 1.195 49.125 1.525 ;
        RECT 48.795 -0.165 49.125 0.165 ;
        RECT 48.8 -8.32 49.12 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.155 10.715 50.485 11.045 ;
        RECT 50.155 9.355 50.485 9.685 ;
        RECT 50.155 7.995 50.485 8.325 ;
        RECT 50.155 6.635 50.485 6.965 ;
        RECT 50.155 5.275 50.485 5.605 ;
        RECT 50.155 3.915 50.485 4.245 ;
        RECT 50.155 2.555 50.485 2.885 ;
        RECT 50.155 1.195 50.485 1.525 ;
        RECT 50.155 -0.165 50.485 0.165 ;
        RECT 50.16 -8.32 50.48 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.515 10.715 51.845 11.045 ;
        RECT 51.515 9.355 51.845 9.685 ;
        RECT 51.515 7.995 51.845 8.325 ;
        RECT 51.515 6.635 51.845 6.965 ;
        RECT 51.515 5.275 51.845 5.605 ;
        RECT 51.515 3.915 51.845 4.245 ;
        RECT 51.515 2.555 51.845 2.885 ;
        RECT 51.515 1.195 51.845 1.525 ;
        RECT 51.515 -0.165 51.845 0.165 ;
        RECT 51.52 -8.32 51.84 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.875 10.715 53.205 11.045 ;
        RECT 52.875 9.355 53.205 9.685 ;
        RECT 52.875 7.995 53.205 8.325 ;
        RECT 52.875 6.635 53.205 6.965 ;
        RECT 52.875 5.275 53.205 5.605 ;
        RECT 52.875 3.915 53.205 4.245 ;
        RECT 52.875 2.555 53.205 2.885 ;
        RECT 52.875 1.195 53.205 1.525 ;
        RECT 52.875 -0.165 53.205 0.165 ;
        RECT 52.88 -8.32 53.2 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.235 10.715 54.565 11.045 ;
        RECT 54.235 9.355 54.565 9.685 ;
        RECT 54.235 7.995 54.565 8.325 ;
        RECT 54.235 6.635 54.565 6.965 ;
        RECT 54.235 5.275 54.565 5.605 ;
        RECT 54.235 3.915 54.565 4.245 ;
        RECT 54.235 2.555 54.565 2.885 ;
        RECT 54.235 1.195 54.565 1.525 ;
        RECT 54.235 -0.165 54.565 0.165 ;
        RECT 54.24 -8.32 54.56 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.595 10.715 55.925 11.045 ;
        RECT 55.595 9.355 55.925 9.685 ;
        RECT 55.595 7.995 55.925 8.325 ;
        RECT 55.595 6.635 55.925 6.965 ;
        RECT 55.595 5.275 55.925 5.605 ;
        RECT 55.595 3.915 55.925 4.245 ;
        RECT 55.595 2.555 55.925 2.885 ;
        RECT 55.595 1.195 55.925 1.525 ;
        RECT 55.595 -0.165 55.925 0.165 ;
        RECT 55.6 -8.32 55.92 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.955 10.715 57.285 11.045 ;
        RECT 56.955 9.355 57.285 9.685 ;
        RECT 56.955 7.995 57.285 8.325 ;
        RECT 56.955 6.635 57.285 6.965 ;
        RECT 56.955 5.275 57.285 5.605 ;
        RECT 56.955 3.915 57.285 4.245 ;
        RECT 56.955 2.555 57.285 2.885 ;
        RECT 56.955 1.195 57.285 1.525 ;
        RECT 56.955 -0.165 57.285 0.165 ;
        RECT 56.96 -8.32 57.28 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.315 10.715 58.645 11.045 ;
        RECT 58.315 9.355 58.645 9.685 ;
        RECT 58.315 7.995 58.645 8.325 ;
        RECT 58.315 6.635 58.645 6.965 ;
        RECT 58.315 5.275 58.645 5.605 ;
        RECT 58.315 3.915 58.645 4.245 ;
        RECT 58.315 2.555 58.645 2.885 ;
        RECT 58.315 1.195 58.645 1.525 ;
        RECT 58.315 -0.165 58.645 0.165 ;
        RECT 58.32 -8.32 58.64 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.675 10.715 60.005 11.045 ;
        RECT 59.675 9.355 60.005 9.685 ;
        RECT 59.675 7.995 60.005 8.325 ;
        RECT 59.675 6.635 60.005 6.965 ;
        RECT 59.675 5.275 60.005 5.605 ;
        RECT 59.675 3.915 60.005 4.245 ;
        RECT 59.675 2.555 60.005 2.885 ;
        RECT 59.675 1.195 60.005 1.525 ;
        RECT 59.675 -0.165 60.005 0.165 ;
        RECT 59.68 -8.32 60 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.035 10.715 61.365 11.045 ;
        RECT 61.035 9.355 61.365 9.685 ;
        RECT 61.035 7.995 61.365 8.325 ;
        RECT 61.035 6.635 61.365 6.965 ;
        RECT 61.035 5.275 61.365 5.605 ;
        RECT 61.035 3.915 61.365 4.245 ;
        RECT 61.035 2.555 61.365 2.885 ;
        RECT 61.035 1.195 61.365 1.525 ;
        RECT 61.035 -0.165 61.365 0.165 ;
        RECT 61.04 -8.32 61.36 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.395 10.715 62.725 11.045 ;
        RECT 62.395 9.355 62.725 9.685 ;
        RECT 62.395 7.995 62.725 8.325 ;
        RECT 62.395 6.635 62.725 6.965 ;
        RECT 62.395 5.275 62.725 5.605 ;
        RECT 62.395 3.915 62.725 4.245 ;
        RECT 62.395 2.555 62.725 2.885 ;
        RECT 62.395 1.195 62.725 1.525 ;
        RECT 62.395 -0.165 62.725 0.165 ;
        RECT 62.4 -8.32 62.72 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.755 10.715 64.085 11.045 ;
        RECT 63.755 9.355 64.085 9.685 ;
        RECT 63.755 7.995 64.085 8.325 ;
        RECT 63.755 6.635 64.085 6.965 ;
        RECT 63.755 5.275 64.085 5.605 ;
        RECT 63.755 3.915 64.085 4.245 ;
        RECT 63.755 2.555 64.085 2.885 ;
        RECT 63.755 1.195 64.085 1.525 ;
        RECT 63.755 -0.165 64.085 0.165 ;
        RECT 63.76 -8.32 64.08 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.115 10.715 65.445 11.045 ;
        RECT 65.115 9.355 65.445 9.685 ;
        RECT 65.115 7.995 65.445 8.325 ;
        RECT 65.115 6.635 65.445 6.965 ;
        RECT 65.115 5.275 65.445 5.605 ;
        RECT 65.115 3.915 65.445 4.245 ;
        RECT 65.115 2.555 65.445 2.885 ;
        RECT 65.115 1.195 65.445 1.525 ;
        RECT 65.115 -0.165 65.445 0.165 ;
        RECT 65.12 -8.32 65.44 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.475 10.715 66.805 11.045 ;
        RECT 66.475 9.355 66.805 9.685 ;
        RECT 66.475 7.995 66.805 8.325 ;
        RECT 66.475 6.635 66.805 6.965 ;
        RECT 66.475 5.275 66.805 5.605 ;
        RECT 66.475 3.915 66.805 4.245 ;
        RECT 66.475 2.555 66.805 2.885 ;
        RECT 66.475 1.195 66.805 1.525 ;
        RECT 66.475 -0.165 66.805 0.165 ;
        RECT 66.48 -8.32 66.8 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.835 10.715 68.165 11.045 ;
        RECT 67.835 9.355 68.165 9.685 ;
        RECT 67.835 7.995 68.165 8.325 ;
        RECT 67.835 6.635 68.165 6.965 ;
        RECT 67.835 5.275 68.165 5.605 ;
        RECT 67.835 3.915 68.165 4.245 ;
        RECT 67.835 2.555 68.165 2.885 ;
        RECT 67.835 1.195 68.165 1.525 ;
        RECT 67.835 -0.165 68.165 0.165 ;
        RECT 67.84 -8.32 68.16 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.195 10.715 69.525 11.045 ;
        RECT 69.195 9.355 69.525 9.685 ;
        RECT 69.195 7.995 69.525 8.325 ;
        RECT 69.195 6.635 69.525 6.965 ;
        RECT 69.195 5.275 69.525 5.605 ;
        RECT 69.195 3.915 69.525 4.245 ;
        RECT 69.195 2.555 69.525 2.885 ;
        RECT 69.195 1.195 69.525 1.525 ;
        RECT 69.195 -0.165 69.525 0.165 ;
        RECT 69.2 -8.32 69.52 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.555 10.715 70.885 11.045 ;
        RECT 70.555 9.355 70.885 9.685 ;
        RECT 70.555 7.995 70.885 8.325 ;
        RECT 70.555 6.635 70.885 6.965 ;
        RECT 70.555 5.275 70.885 5.605 ;
        RECT 70.555 3.915 70.885 4.245 ;
        RECT 70.555 2.555 70.885 2.885 ;
        RECT 70.555 1.195 70.885 1.525 ;
        RECT 70.555 -0.165 70.885 0.165 ;
        RECT 70.56 -8.32 70.88 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915 10.715 72.245 11.045 ;
        RECT 71.915 9.355 72.245 9.685 ;
        RECT 71.915 7.995 72.245 8.325 ;
        RECT 71.915 6.635 72.245 6.965 ;
        RECT 71.915 5.275 72.245 5.605 ;
        RECT 71.915 3.915 72.245 4.245 ;
        RECT 71.915 2.555 72.245 2.885 ;
        RECT 71.915 1.195 72.245 1.525 ;
        RECT 71.915 -0.165 72.245 0.165 ;
        RECT 71.92 -8.32 72.24 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.275 10.715 73.605 11.045 ;
        RECT 73.275 9.355 73.605 9.685 ;
        RECT 73.275 7.995 73.605 8.325 ;
        RECT 73.275 6.635 73.605 6.965 ;
        RECT 73.275 5.275 73.605 5.605 ;
        RECT 73.275 3.915 73.605 4.245 ;
        RECT 73.275 2.555 73.605 2.885 ;
        RECT 73.275 1.195 73.605 1.525 ;
        RECT 73.275 -0.165 73.605 0.165 ;
        RECT 73.28 -8.32 73.6 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.635 10.715 74.965 11.045 ;
        RECT 74.635 9.355 74.965 9.685 ;
        RECT 74.635 7.995 74.965 8.325 ;
        RECT 74.635 6.635 74.965 6.965 ;
        RECT 74.635 5.275 74.965 5.605 ;
        RECT 74.635 3.915 74.965 4.245 ;
        RECT 74.635 2.555 74.965 2.885 ;
        RECT 74.635 1.195 74.965 1.525 ;
        RECT 74.635 -0.165 74.965 0.165 ;
        RECT 74.64 -8.32 74.96 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.995 10.715 76.325 11.045 ;
        RECT 75.995 9.355 76.325 9.685 ;
        RECT 75.995 7.995 76.325 8.325 ;
        RECT 75.995 6.635 76.325 6.965 ;
        RECT 75.995 5.275 76.325 5.605 ;
        RECT 75.995 3.915 76.325 4.245 ;
        RECT 75.995 2.555 76.325 2.885 ;
        RECT 75.995 1.195 76.325 1.525 ;
        RECT 75.995 -0.165 76.325 0.165 ;
        RECT 76 -8.32 76.32 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.355 10.715 77.685 11.045 ;
        RECT 77.355 9.355 77.685 9.685 ;
        RECT 77.355 7.995 77.685 8.325 ;
        RECT 77.355 6.635 77.685 6.965 ;
        RECT 77.355 5.275 77.685 5.605 ;
        RECT 77.355 3.915 77.685 4.245 ;
        RECT 77.355 2.555 77.685 2.885 ;
        RECT 77.355 1.195 77.685 1.525 ;
        RECT 77.355 -0.165 77.685 0.165 ;
        RECT 77.36 -8.32 77.68 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.715 10.715 79.045 11.045 ;
        RECT 78.715 9.355 79.045 9.685 ;
        RECT 78.715 7.995 79.045 8.325 ;
        RECT 78.715 6.635 79.045 6.965 ;
        RECT 78.715 5.275 79.045 5.605 ;
        RECT 78.715 3.915 79.045 4.245 ;
        RECT 78.715 2.555 79.045 2.885 ;
        RECT 78.715 1.195 79.045 1.525 ;
        RECT 78.715 -0.165 79.045 0.165 ;
        RECT 78.72 -8.32 79.04 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.075 10.715 80.405 11.045 ;
        RECT 80.075 9.355 80.405 9.685 ;
        RECT 80.075 7.995 80.405 8.325 ;
        RECT 80.075 6.635 80.405 6.965 ;
        RECT 80.075 5.275 80.405 5.605 ;
        RECT 80.075 3.915 80.405 4.245 ;
        RECT 80.075 2.555 80.405 2.885 ;
        RECT 80.075 1.195 80.405 1.525 ;
        RECT 80.075 -0.165 80.405 0.165 ;
        RECT 80.08 -8.32 80.4 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.435 10.715 81.765 11.045 ;
        RECT 81.435 9.355 81.765 9.685 ;
        RECT 81.435 7.995 81.765 8.325 ;
        RECT 81.435 6.635 81.765 6.965 ;
        RECT 81.435 5.275 81.765 5.605 ;
        RECT 81.435 3.915 81.765 4.245 ;
        RECT 81.435 2.555 81.765 2.885 ;
        RECT 81.435 1.195 81.765 1.525 ;
        RECT 81.435 -0.165 81.765 0.165 ;
        RECT 81.44 -8.32 81.76 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.795 10.715 83.125 11.045 ;
        RECT 82.795 9.355 83.125 9.685 ;
        RECT 82.795 7.995 83.125 8.325 ;
        RECT 82.795 6.635 83.125 6.965 ;
        RECT 82.795 5.275 83.125 5.605 ;
        RECT 82.795 3.915 83.125 4.245 ;
        RECT 82.795 2.555 83.125 2.885 ;
        RECT 82.795 1.195 83.125 1.525 ;
        RECT 82.795 -0.165 83.125 0.165 ;
        RECT 82.8 -8.32 83.12 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.155 10.715 84.485 11.045 ;
        RECT 84.155 9.355 84.485 9.685 ;
        RECT 84.155 7.995 84.485 8.325 ;
        RECT 84.155 6.635 84.485 6.965 ;
        RECT 84.155 5.275 84.485 5.605 ;
        RECT 84.155 3.915 84.485 4.245 ;
        RECT 84.155 2.555 84.485 2.885 ;
        RECT 84.155 1.195 84.485 1.525 ;
        RECT 84.155 -0.165 84.485 0.165 ;
        RECT 84.16 -8.32 84.48 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.515 10.715 85.845 11.045 ;
        RECT 85.515 9.355 85.845 9.685 ;
        RECT 85.515 7.995 85.845 8.325 ;
        RECT 85.515 6.635 85.845 6.965 ;
        RECT 85.515 5.275 85.845 5.605 ;
        RECT 85.515 3.915 85.845 4.245 ;
        RECT 85.515 2.555 85.845 2.885 ;
        RECT 85.515 1.195 85.845 1.525 ;
        RECT 85.515 -0.165 85.845 0.165 ;
        RECT 85.52 -8.32 85.84 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.875 10.715 87.205 11.045 ;
        RECT 86.875 9.355 87.205 9.685 ;
        RECT 86.875 7.995 87.205 8.325 ;
        RECT 86.875 6.635 87.205 6.965 ;
        RECT 86.875 5.275 87.205 5.605 ;
        RECT 86.875 3.915 87.205 4.245 ;
        RECT 86.875 2.555 87.205 2.885 ;
        RECT 86.875 1.195 87.205 1.525 ;
        RECT 86.875 -0.165 87.205 0.165 ;
        RECT 86.88 -8.32 87.2 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.235 10.715 88.565 11.045 ;
        RECT 88.235 9.355 88.565 9.685 ;
        RECT 88.235 7.995 88.565 8.325 ;
        RECT 88.235 6.635 88.565 6.965 ;
        RECT 88.235 5.275 88.565 5.605 ;
        RECT 88.235 3.915 88.565 4.245 ;
        RECT 88.235 2.555 88.565 2.885 ;
        RECT 88.235 1.195 88.565 1.525 ;
        RECT 88.235 -0.165 88.565 0.165 ;
        RECT 88.24 -8.32 88.56 15.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 89.595 9.355 89.925 9.685 ;
        RECT 89.595 7.995 89.925 8.325 ;
        RECT 89.595 6.635 89.925 6.965 ;
        RECT 89.595 5.275 89.925 5.605 ;
        RECT 89.595 3.915 89.925 4.245 ;
        RECT 89.595 2.555 89.925 2.885 ;
        RECT 89.595 1.195 89.925 1.525 ;
        RECT 89.595 -0.165 89.925 0.165 ;
        RECT 89.6 -8.32 89.92 15.8 ;
        RECT 89.595 10.715 89.925 11.045 ;
    END
  END vss
  OBS
    LAYER met1 SPACING 0.14 ;
      RECT 0.88 0 766.87 6.92 ;
    LAYER met2 SPACING 0.14 ;
      RECT -2.91 -8.32 769.27 15.8 ;
  END
END tristate_inv_delay_line_128

END LIBRARY
