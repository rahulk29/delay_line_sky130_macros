VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO tristate_inv_delay_line_128
  CLASS BLOCK ;
  ORIGIN 2.225 1.525 ;
  FOREIGN tristate_inv_delay_line_128 -2.225 -1.525 ;
  SIZE 771.49 BY 10.53 ;
  SYMMETRY X Y R90 ;
  PIN clk_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT -0.47 0 -0.15 0.32 ;
    END
  END clk_in
  PIN clk_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.52 0 1.84 0.32 ;
    END
  END clk_out
  PIN ctl[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.03 0 0.35 0.32 ;
    END
  END ctl[0]
  PIN ctl[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 600.03 0 600.35 0.32 ;
    END
  END ctl[100]
  PIN ctl[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 606.03 0 606.35 0.32 ;
    END
  END ctl[101]
  PIN ctl[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 612.03 0 612.35 0.32 ;
    END
  END ctl[102]
  PIN ctl[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 618.03 0 618.35 0.32 ;
    END
  END ctl[103]
  PIN ctl[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 624.03 0 624.35 0.32 ;
    END
  END ctl[104]
  PIN ctl[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 630.03 0 630.35 0.32 ;
    END
  END ctl[105]
  PIN ctl[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 636.03 0 636.35 0.32 ;
    END
  END ctl[106]
  PIN ctl[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 642.03 0 642.35 0.32 ;
    END
  END ctl[107]
  PIN ctl[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 648.03 0 648.35 0.32 ;
    END
  END ctl[108]
  PIN ctl[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 654.03 0 654.35 0.32 ;
    END
  END ctl[109]
  PIN ctl[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 60.03 0 60.35 0.32 ;
    END
  END ctl[10]
  PIN ctl[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 660.03 0 660.35 0.32 ;
    END
  END ctl[110]
  PIN ctl[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 666.03 0 666.35 0.32 ;
    END
  END ctl[111]
  PIN ctl[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 672.03 0 672.35 0.32 ;
    END
  END ctl[112]
  PIN ctl[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 678.03 0 678.35 0.32 ;
    END
  END ctl[113]
  PIN ctl[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 684.03 0 684.35 0.32 ;
    END
  END ctl[114]
  PIN ctl[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 690.03 0 690.35 0.32 ;
    END
  END ctl[115]
  PIN ctl[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 696.03 0 696.35 0.32 ;
    END
  END ctl[116]
  PIN ctl[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 702.03 0 702.35 0.32 ;
    END
  END ctl[117]
  PIN ctl[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 708.03 0 708.35 0.32 ;
    END
  END ctl[118]
  PIN ctl[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 714.03 0 714.35 0.32 ;
    END
  END ctl[119]
  PIN ctl[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 66.03 0 66.35 0.32 ;
    END
  END ctl[11]
  PIN ctl[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 720.03 0 720.35 0.32 ;
    END
  END ctl[120]
  PIN ctl[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 726.03 0 726.35 0.32 ;
    END
  END ctl[121]
  PIN ctl[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 732.03 0 732.35 0.32 ;
    END
  END ctl[122]
  PIN ctl[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 738.03 0 738.35 0.32 ;
    END
  END ctl[123]
  PIN ctl[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 744.03 0 744.35 0.32 ;
    END
  END ctl[124]
  PIN ctl[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 750.03 0 750.35 0.32 ;
    END
  END ctl[125]
  PIN ctl[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 756.03 0 756.35 0.32 ;
    END
  END ctl[126]
  PIN ctl[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 762.03 0 762.35 0.32 ;
    END
  END ctl[127]
  PIN ctl[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 72.03 0 72.35 0.32 ;
    END
  END ctl[12]
  PIN ctl[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 78.03 0 78.35 0.32 ;
    END
  END ctl[13]
  PIN ctl[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 84.03 0 84.35 0.32 ;
    END
  END ctl[14]
  PIN ctl[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 90.03 0 90.35 0.32 ;
    END
  END ctl[15]
  PIN ctl[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 96.03 0 96.35 0.32 ;
    END
  END ctl[16]
  PIN ctl[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 102.03 0 102.35 0.32 ;
    END
  END ctl[17]
  PIN ctl[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 108.03 0 108.35 0.32 ;
    END
  END ctl[18]
  PIN ctl[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 114.03 0 114.35 0.32 ;
    END
  END ctl[19]
  PIN ctl[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 6.03 0 6.35 0.32 ;
    END
  END ctl[1]
  PIN ctl[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 120.03 0 120.35 0.32 ;
    END
  END ctl[20]
  PIN ctl[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 126.03 0 126.35 0.32 ;
    END
  END ctl[21]
  PIN ctl[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 132.03 0 132.35 0.32 ;
    END
  END ctl[22]
  PIN ctl[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 138.03 0 138.35 0.32 ;
    END
  END ctl[23]
  PIN ctl[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 144.03 0 144.35 0.32 ;
    END
  END ctl[24]
  PIN ctl[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 150.03 0 150.35 0.32 ;
    END
  END ctl[25]
  PIN ctl[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 156.03 0 156.35 0.32 ;
    END
  END ctl[26]
  PIN ctl[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 162.03 0 162.35 0.32 ;
    END
  END ctl[27]
  PIN ctl[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 168.03 0 168.35 0.32 ;
    END
  END ctl[28]
  PIN ctl[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 174.03 0 174.35 0.32 ;
    END
  END ctl[29]
  PIN ctl[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 12.03 0 12.35 0.32 ;
    END
  END ctl[2]
  PIN ctl[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 180.03 0 180.35 0.32 ;
    END
  END ctl[30]
  PIN ctl[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 186.03 0 186.35 0.32 ;
    END
  END ctl[31]
  PIN ctl[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 192.03 0 192.35 0.32 ;
    END
  END ctl[32]
  PIN ctl[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 198.03 0 198.35 0.32 ;
    END
  END ctl[33]
  PIN ctl[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 204.03 0 204.35 0.32 ;
    END
  END ctl[34]
  PIN ctl[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 210.03 0 210.35 0.32 ;
    END
  END ctl[35]
  PIN ctl[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 216.03 0 216.35 0.32 ;
    END
  END ctl[36]
  PIN ctl[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 222.03 0 222.35 0.32 ;
    END
  END ctl[37]
  PIN ctl[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 228.03 0 228.35 0.32 ;
    END
  END ctl[38]
  PIN ctl[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 234.03 0 234.35 0.32 ;
    END
  END ctl[39]
  PIN ctl[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.03 0 18.35 0.32 ;
    END
  END ctl[3]
  PIN ctl[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 240.03 0 240.35 0.32 ;
    END
  END ctl[40]
  PIN ctl[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 246.03 0 246.35 0.32 ;
    END
  END ctl[41]
  PIN ctl[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 252.03 0 252.35 0.32 ;
    END
  END ctl[42]
  PIN ctl[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 258.03 0 258.35 0.32 ;
    END
  END ctl[43]
  PIN ctl[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 264.03 0 264.35 0.32 ;
    END
  END ctl[44]
  PIN ctl[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 270.03 0 270.35 0.32 ;
    END
  END ctl[45]
  PIN ctl[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 276.03 0 276.35 0.32 ;
    END
  END ctl[46]
  PIN ctl[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 282.03 0 282.35 0.32 ;
    END
  END ctl[47]
  PIN ctl[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 288.03 0 288.35 0.32 ;
    END
  END ctl[48]
  PIN ctl[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 294.03 0 294.35 0.32 ;
    END
  END ctl[49]
  PIN ctl[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 24.03 0 24.35 0.32 ;
    END
  END ctl[4]
  PIN ctl[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 300.03 0 300.35 0.32 ;
    END
  END ctl[50]
  PIN ctl[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 306.03 0 306.35 0.32 ;
    END
  END ctl[51]
  PIN ctl[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 312.03 0 312.35 0.32 ;
    END
  END ctl[52]
  PIN ctl[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 318.03 0 318.35 0.32 ;
    END
  END ctl[53]
  PIN ctl[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 324.03 0 324.35 0.32 ;
    END
  END ctl[54]
  PIN ctl[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 330.03 0 330.35 0.32 ;
    END
  END ctl[55]
  PIN ctl[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 336.03 0 336.35 0.32 ;
    END
  END ctl[56]
  PIN ctl[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 342.03 0 342.35 0.32 ;
    END
  END ctl[57]
  PIN ctl[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 348.03 0 348.35 0.32 ;
    END
  END ctl[58]
  PIN ctl[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 354.03 0 354.35 0.32 ;
    END
  END ctl[59]
  PIN ctl[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 30.03 0 30.35 0.32 ;
    END
  END ctl[5]
  PIN ctl[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 360.03 0 360.35 0.32 ;
    END
  END ctl[60]
  PIN ctl[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 366.03 0 366.35 0.32 ;
    END
  END ctl[61]
  PIN ctl[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 372.03 0 372.35 0.32 ;
    END
  END ctl[62]
  PIN ctl[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 378.03 0 378.35 0.32 ;
    END
  END ctl[63]
  PIN ctl[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 384.03 0 384.35 0.32 ;
    END
  END ctl[64]
  PIN ctl[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 390.03 0 390.35 0.32 ;
    END
  END ctl[65]
  PIN ctl[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 396.03 0 396.35 0.32 ;
    END
  END ctl[66]
  PIN ctl[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 402.03 0 402.35 0.32 ;
    END
  END ctl[67]
  PIN ctl[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 408.03 0 408.35 0.32 ;
    END
  END ctl[68]
  PIN ctl[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 414.03 0 414.35 0.32 ;
    END
  END ctl[69]
  PIN ctl[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 36.03 0 36.35 0.32 ;
    END
  END ctl[6]
  PIN ctl[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 420.03 0 420.35 0.32 ;
    END
  END ctl[70]
  PIN ctl[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 426.03 0 426.35 0.32 ;
    END
  END ctl[71]
  PIN ctl[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 432.03 0 432.35 0.32 ;
    END
  END ctl[72]
  PIN ctl[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 438.03 0 438.35 0.32 ;
    END
  END ctl[73]
  PIN ctl[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 444.03 0 444.35 0.32 ;
    END
  END ctl[74]
  PIN ctl[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 450.03 0 450.35 0.32 ;
    END
  END ctl[75]
  PIN ctl[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 456.03 0 456.35 0.32 ;
    END
  END ctl[76]
  PIN ctl[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 462.03 0 462.35 0.32 ;
    END
  END ctl[77]
  PIN ctl[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 468.03 0 468.35 0.32 ;
    END
  END ctl[78]
  PIN ctl[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 474.03 0 474.35 0.32 ;
    END
  END ctl[79]
  PIN ctl[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 42.03 0 42.35 0.32 ;
    END
  END ctl[7]
  PIN ctl[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 480.03 0 480.35 0.32 ;
    END
  END ctl[80]
  PIN ctl[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 486.03 0 486.35 0.32 ;
    END
  END ctl[81]
  PIN ctl[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 492.03 0 492.35 0.32 ;
    END
  END ctl[82]
  PIN ctl[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 498.03 0 498.35 0.32 ;
    END
  END ctl[83]
  PIN ctl[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 504.03 0 504.35 0.32 ;
    END
  END ctl[84]
  PIN ctl[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 510.03 0 510.35 0.32 ;
    END
  END ctl[85]
  PIN ctl[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 516.03 0 516.35 0.32 ;
    END
  END ctl[86]
  PIN ctl[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 522.03 0 522.35 0.32 ;
    END
  END ctl[87]
  PIN ctl[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 528.03 0 528.35 0.32 ;
    END
  END ctl[88]
  PIN ctl[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 534.03 0 534.35 0.32 ;
    END
  END ctl[89]
  PIN ctl[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 48.03 0 48.35 0.32 ;
    END
  END ctl[8]
  PIN ctl[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 540.03 0 540.35 0.32 ;
    END
  END ctl[90]
  PIN ctl[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 546.03 0 546.35 0.32 ;
    END
  END ctl[91]
  PIN ctl[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 552.03 0 552.35 0.32 ;
    END
  END ctl[92]
  PIN ctl[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 558.03 0 558.35 0.32 ;
    END
  END ctl[93]
  PIN ctl[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 564.03 0 564.35 0.32 ;
    END
  END ctl[94]
  PIN ctl[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 570.03 0 570.35 0.32 ;
    END
  END ctl[95]
  PIN ctl[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 576.03 0 576.35 0.32 ;
    END
  END ctl[96]
  PIN ctl[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 582.03 0 582.35 0.32 ;
    END
  END ctl[97]
  PIN ctl[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 588.03 0 588.35 0.32 ;
    END
  END ctl[98]
  PIN ctl[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 594.03 0 594.35 0.32 ;
    END
  END ctl[99]
  PIN ctl[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 54.03 0 54.35 0.32 ;
    END
  END ctl[9]
  PIN ctl_b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 4.05 0 4.37 0.32 ;
    END
  END ctl_b[0]
  PIN ctl_b[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 604.05 0 604.37 0.32 ;
    END
  END ctl_b[100]
  PIN ctl_b[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 610.05 0 610.37 0.32 ;
    END
  END ctl_b[101]
  PIN ctl_b[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 616.05 0 616.37 0.32 ;
    END
  END ctl_b[102]
  PIN ctl_b[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 622.05 0 622.37 0.32 ;
    END
  END ctl_b[103]
  PIN ctl_b[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 628.05 0 628.37 0.32 ;
    END
  END ctl_b[104]
  PIN ctl_b[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 634.05 0 634.37 0.32 ;
    END
  END ctl_b[105]
  PIN ctl_b[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 640.05 0 640.37 0.32 ;
    END
  END ctl_b[106]
  PIN ctl_b[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 646.05 0 646.37 0.32 ;
    END
  END ctl_b[107]
  PIN ctl_b[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 652.05 0 652.37 0.32 ;
    END
  END ctl_b[108]
  PIN ctl_b[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 658.05 0 658.37 0.32 ;
    END
  END ctl_b[109]
  PIN ctl_b[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 64.05 0 64.37 0.32 ;
    END
  END ctl_b[10]
  PIN ctl_b[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 664.05 0 664.37 0.32 ;
    END
  END ctl_b[110]
  PIN ctl_b[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 670.05 0 670.37 0.32 ;
    END
  END ctl_b[111]
  PIN ctl_b[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 676.05 0 676.37 0.32 ;
    END
  END ctl_b[112]
  PIN ctl_b[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 682.05 0 682.37 0.32 ;
    END
  END ctl_b[113]
  PIN ctl_b[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 688.05 0 688.37 0.32 ;
    END
  END ctl_b[114]
  PIN ctl_b[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 694.05 0 694.37 0.32 ;
    END
  END ctl_b[115]
  PIN ctl_b[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 700.05 0 700.37 0.32 ;
    END
  END ctl_b[116]
  PIN ctl_b[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 706.05 0 706.37 0.32 ;
    END
  END ctl_b[117]
  PIN ctl_b[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 712.05 0 712.37 0.32 ;
    END
  END ctl_b[118]
  PIN ctl_b[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 718.05 0 718.37 0.32 ;
    END
  END ctl_b[119]
  PIN ctl_b[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 70.05 0 70.37 0.32 ;
    END
  END ctl_b[11]
  PIN ctl_b[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 724.05 0 724.37 0.32 ;
    END
  END ctl_b[120]
  PIN ctl_b[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 730.05 0 730.37 0.32 ;
    END
  END ctl_b[121]
  PIN ctl_b[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 736.05 0 736.37 0.32 ;
    END
  END ctl_b[122]
  PIN ctl_b[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 742.05 0 742.37 0.32 ;
    END
  END ctl_b[123]
  PIN ctl_b[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 748.05 0 748.37 0.32 ;
    END
  END ctl_b[124]
  PIN ctl_b[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 754.05 0 754.37 0.32 ;
    END
  END ctl_b[125]
  PIN ctl_b[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 760.05 0 760.37 0.32 ;
    END
  END ctl_b[126]
  PIN ctl_b[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 766.05 0 766.37 0.32 ;
    END
  END ctl_b[127]
  PIN ctl_b[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 76.05 0 76.37 0.32 ;
    END
  END ctl_b[12]
  PIN ctl_b[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 82.05 0 82.37 0.32 ;
    END
  END ctl_b[13]
  PIN ctl_b[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 88.05 0 88.37 0.32 ;
    END
  END ctl_b[14]
  PIN ctl_b[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 94.05 0 94.37 0.32 ;
    END
  END ctl_b[15]
  PIN ctl_b[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 100.05 0 100.37 0.32 ;
    END
  END ctl_b[16]
  PIN ctl_b[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 106.05 0 106.37 0.32 ;
    END
  END ctl_b[17]
  PIN ctl_b[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 112.05 0 112.37 0.32 ;
    END
  END ctl_b[18]
  PIN ctl_b[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 118.05 0 118.37 0.32 ;
    END
  END ctl_b[19]
  PIN ctl_b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 10.05 0 10.37 0.32 ;
    END
  END ctl_b[1]
  PIN ctl_b[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 124.05 0 124.37 0.32 ;
    END
  END ctl_b[20]
  PIN ctl_b[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 130.05 0 130.37 0.32 ;
    END
  END ctl_b[21]
  PIN ctl_b[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 136.05 0 136.37 0.32 ;
    END
  END ctl_b[22]
  PIN ctl_b[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 142.05 0 142.37 0.32 ;
    END
  END ctl_b[23]
  PIN ctl_b[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 148.05 0 148.37 0.32 ;
    END
  END ctl_b[24]
  PIN ctl_b[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 154.05 0 154.37 0.32 ;
    END
  END ctl_b[25]
  PIN ctl_b[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 160.05 0 160.37 0.32 ;
    END
  END ctl_b[26]
  PIN ctl_b[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 166.05 0 166.37 0.32 ;
    END
  END ctl_b[27]
  PIN ctl_b[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 172.05 0 172.37 0.32 ;
    END
  END ctl_b[28]
  PIN ctl_b[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 178.05 0 178.37 0.32 ;
    END
  END ctl_b[29]
  PIN ctl_b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.05 0 16.37 0.32 ;
    END
  END ctl_b[2]
  PIN ctl_b[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 184.05 0 184.37 0.32 ;
    END
  END ctl_b[30]
  PIN ctl_b[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 190.05 0 190.37 0.32 ;
    END
  END ctl_b[31]
  PIN ctl_b[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 196.05 0 196.37 0.32 ;
    END
  END ctl_b[32]
  PIN ctl_b[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 202.05 0 202.37 0.32 ;
    END
  END ctl_b[33]
  PIN ctl_b[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 208.05 0 208.37 0.32 ;
    END
  END ctl_b[34]
  PIN ctl_b[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 214.05 0 214.37 0.32 ;
    END
  END ctl_b[35]
  PIN ctl_b[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 220.05 0 220.37 0.32 ;
    END
  END ctl_b[36]
  PIN ctl_b[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 226.05 0 226.37 0.32 ;
    END
  END ctl_b[37]
  PIN ctl_b[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 232.05 0 232.37 0.32 ;
    END
  END ctl_b[38]
  PIN ctl_b[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 238.05 0 238.37 0.32 ;
    END
  END ctl_b[39]
  PIN ctl_b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 22.05 0 22.37 0.32 ;
    END
  END ctl_b[3]
  PIN ctl_b[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 244.05 0 244.37 0.32 ;
    END
  END ctl_b[40]
  PIN ctl_b[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 250.05 0 250.37 0.32 ;
    END
  END ctl_b[41]
  PIN ctl_b[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 256.05 0 256.37 0.32 ;
    END
  END ctl_b[42]
  PIN ctl_b[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 262.05 0 262.37 0.32 ;
    END
  END ctl_b[43]
  PIN ctl_b[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 268.05 0 268.37 0.32 ;
    END
  END ctl_b[44]
  PIN ctl_b[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 274.05 0 274.37 0.32 ;
    END
  END ctl_b[45]
  PIN ctl_b[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 280.05 0 280.37 0.32 ;
    END
  END ctl_b[46]
  PIN ctl_b[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 286.05 0 286.37 0.32 ;
    END
  END ctl_b[47]
  PIN ctl_b[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 292.05 0 292.37 0.32 ;
    END
  END ctl_b[48]
  PIN ctl_b[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 298.05 0 298.37 0.32 ;
    END
  END ctl_b[49]
  PIN ctl_b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 28.05 0 28.37 0.32 ;
    END
  END ctl_b[4]
  PIN ctl_b[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 304.05 0 304.37 0.32 ;
    END
  END ctl_b[50]
  PIN ctl_b[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 310.05 0 310.37 0.32 ;
    END
  END ctl_b[51]
  PIN ctl_b[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 316.05 0 316.37 0.32 ;
    END
  END ctl_b[52]
  PIN ctl_b[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 322.05 0 322.37 0.32 ;
    END
  END ctl_b[53]
  PIN ctl_b[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 328.05 0 328.37 0.32 ;
    END
  END ctl_b[54]
  PIN ctl_b[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 334.05 0 334.37 0.32 ;
    END
  END ctl_b[55]
  PIN ctl_b[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 340.05 0 340.37 0.32 ;
    END
  END ctl_b[56]
  PIN ctl_b[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 346.05 0 346.37 0.32 ;
    END
  END ctl_b[57]
  PIN ctl_b[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 352.05 0 352.37 0.32 ;
    END
  END ctl_b[58]
  PIN ctl_b[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 358.05 0 358.37 0.32 ;
    END
  END ctl_b[59]
  PIN ctl_b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 34.05 0 34.37 0.32 ;
    END
  END ctl_b[5]
  PIN ctl_b[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 364.05 0 364.37 0.32 ;
    END
  END ctl_b[60]
  PIN ctl_b[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 370.05 0 370.37 0.32 ;
    END
  END ctl_b[61]
  PIN ctl_b[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 376.05 0 376.37 0.32 ;
    END
  END ctl_b[62]
  PIN ctl_b[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 382.05 0 382.37 0.32 ;
    END
  END ctl_b[63]
  PIN ctl_b[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 388.05 0 388.37 0.32 ;
    END
  END ctl_b[64]
  PIN ctl_b[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 394.05 0 394.37 0.32 ;
    END
  END ctl_b[65]
  PIN ctl_b[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 400.05 0 400.37 0.32 ;
    END
  END ctl_b[66]
  PIN ctl_b[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 406.05 0 406.37 0.32 ;
    END
  END ctl_b[67]
  PIN ctl_b[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 412.05 0 412.37 0.32 ;
    END
  END ctl_b[68]
  PIN ctl_b[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 418.05 0 418.37 0.32 ;
    END
  END ctl_b[69]
  PIN ctl_b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 40.05 0 40.37 0.32 ;
    END
  END ctl_b[6]
  PIN ctl_b[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 424.05 0 424.37 0.32 ;
    END
  END ctl_b[70]
  PIN ctl_b[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 430.05 0 430.37 0.32 ;
    END
  END ctl_b[71]
  PIN ctl_b[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 436.05 0 436.37 0.32 ;
    END
  END ctl_b[72]
  PIN ctl_b[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 442.05 0 442.37 0.32 ;
    END
  END ctl_b[73]
  PIN ctl_b[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 448.05 0 448.37 0.32 ;
    END
  END ctl_b[74]
  PIN ctl_b[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 454.05 0 454.37 0.32 ;
    END
  END ctl_b[75]
  PIN ctl_b[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 460.05 0 460.37 0.32 ;
    END
  END ctl_b[76]
  PIN ctl_b[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 466.05 0 466.37 0.32 ;
    END
  END ctl_b[77]
  PIN ctl_b[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 472.05 0 472.37 0.32 ;
    END
  END ctl_b[78]
  PIN ctl_b[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 478.05 0 478.37 0.32 ;
    END
  END ctl_b[79]
  PIN ctl_b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 46.05 0 46.37 0.32 ;
    END
  END ctl_b[7]
  PIN ctl_b[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 484.05 0 484.37 0.32 ;
    END
  END ctl_b[80]
  PIN ctl_b[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 490.05 0 490.37 0.32 ;
    END
  END ctl_b[81]
  PIN ctl_b[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 496.05 0 496.37 0.32 ;
    END
  END ctl_b[82]
  PIN ctl_b[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 502.05 0 502.37 0.32 ;
    END
  END ctl_b[83]
  PIN ctl_b[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 508.05 0 508.37 0.32 ;
    END
  END ctl_b[84]
  PIN ctl_b[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 514.05 0 514.37 0.32 ;
    END
  END ctl_b[85]
  PIN ctl_b[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 520.05 0 520.37 0.32 ;
    END
  END ctl_b[86]
  PIN ctl_b[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 526.05 0 526.37 0.32 ;
    END
  END ctl_b[87]
  PIN ctl_b[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 532.05 0 532.37 0.32 ;
    END
  END ctl_b[88]
  PIN ctl_b[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 538.05 0 538.37 0.32 ;
    END
  END ctl_b[89]
  PIN ctl_b[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 52.05 0 52.37 0.32 ;
    END
  END ctl_b[8]
  PIN ctl_b[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 544.05 0 544.37 0.32 ;
    END
  END ctl_b[90]
  PIN ctl_b[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 550.05 0 550.37 0.32 ;
    END
  END ctl_b[91]
  PIN ctl_b[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 556.05 0 556.37 0.32 ;
    END
  END ctl_b[92]
  PIN ctl_b[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 562.05 0 562.37 0.32 ;
    END
  END ctl_b[93]
  PIN ctl_b[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 568.05 0 568.37 0.32 ;
    END
  END ctl_b[94]
  PIN ctl_b[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 574.05 0 574.37 0.32 ;
    END
  END ctl_b[95]
  PIN ctl_b[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 580.05 0 580.37 0.32 ;
    END
  END ctl_b[96]
  PIN ctl_b[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 586.05 0 586.37 0.32 ;
    END
  END ctl_b[97]
  PIN ctl_b[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 592.05 0 592.37 0.32 ;
    END
  END ctl_b[98]
  PIN ctl_b[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 598.05 0 598.37 0.32 ;
    END
  END ctl_b[99]
  PIN ctl_b[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 58.05 0 58.37 0.32 ;
    END
  END ctl_b[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 557.435 8.675 557.765 9.005 ;
        RECT 557.435 7.315 557.765 7.645 ;
        RECT 557.435 3.235 557.765 3.565 ;
        RECT 557.435 1.875 557.765 2.205 ;
        RECT 557.435 0.515 557.765 0.845 ;
        RECT 557.435 -0.845 557.765 -0.515 ;
        RECT 557.44 -1.52 557.76 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 558.795 8.675 559.125 9.005 ;
        RECT 558.795 7.315 559.125 7.645 ;
        RECT 558.795 3.235 559.125 3.565 ;
        RECT 558.795 1.875 559.125 2.205 ;
        RECT 558.795 0.515 559.125 0.845 ;
        RECT 558.795 -0.845 559.125 -0.515 ;
        RECT 558.8 -1.52 559.12 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 560.155 8.675 560.485 9.005 ;
        RECT 560.155 7.315 560.485 7.645 ;
        RECT 560.155 1.875 560.485 2.205 ;
        RECT 560.155 0.515 560.485 0.845 ;
        RECT 560.155 -0.845 560.485 -0.515 ;
        RECT 560.16 -1.52 560.48 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 561.515 8.675 561.845 9.005 ;
        RECT 561.515 7.315 561.845 7.645 ;
        RECT 561.515 1.875 561.845 2.205 ;
        RECT 561.515 0.515 561.845 0.845 ;
        RECT 561.515 -0.845 561.845 -0.515 ;
        RECT 561.52 -1.52 561.84 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 562.875 8.675 563.205 9.005 ;
        RECT 562.875 7.315 563.205 7.645 ;
        RECT 562.875 1.875 563.205 2.205 ;
        RECT 562.875 0.515 563.205 0.845 ;
        RECT 562.875 -0.845 563.205 -0.515 ;
        RECT 562.88 -1.52 563.2 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 564.235 8.675 564.565 9.005 ;
        RECT 564.235 7.315 564.565 7.645 ;
        RECT 564.235 1.875 564.565 2.205 ;
        RECT 564.235 0.515 564.565 0.845 ;
        RECT 564.235 -0.845 564.565 -0.515 ;
        RECT 564.24 -1.52 564.56 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 565.595 8.675 565.925 9.005 ;
        RECT 565.595 7.315 565.925 7.645 ;
        RECT 565.595 1.875 565.925 2.205 ;
        RECT 565.595 0.515 565.925 0.845 ;
        RECT 565.595 -0.845 565.925 -0.515 ;
        RECT 565.6 -1.52 565.92 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 566.955 8.675 567.285 9.005 ;
        RECT 566.955 7.315 567.285 7.645 ;
        RECT 566.955 3.235 567.285 3.565 ;
        RECT 566.955 1.875 567.285 2.205 ;
        RECT 566.955 0.515 567.285 0.845 ;
        RECT 566.955 -0.845 567.285 -0.515 ;
        RECT 566.96 -1.52 567.28 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 568.315 8.675 568.645 9.005 ;
        RECT 568.315 7.315 568.645 7.645 ;
        RECT 568.315 3.235 568.645 3.565 ;
        RECT 568.315 1.875 568.645 2.205 ;
        RECT 568.315 0.515 568.645 0.845 ;
        RECT 568.315 -0.845 568.645 -0.515 ;
        RECT 568.32 -1.52 568.64 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 569.675 8.675 570.005 9.005 ;
        RECT 569.675 7.315 570.005 7.645 ;
        RECT 569.675 3.235 570.005 3.565 ;
        RECT 569.675 1.875 570.005 2.205 ;
        RECT 569.675 0.515 570.005 0.845 ;
        RECT 569.675 -0.845 570.005 -0.515 ;
        RECT 569.68 -1.52 570 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 571.035 8.675 571.365 9.005 ;
        RECT 571.035 7.315 571.365 7.645 ;
        RECT 571.035 1.875 571.365 2.205 ;
        RECT 571.035 0.515 571.365 0.845 ;
        RECT 571.035 -0.845 571.365 -0.515 ;
        RECT 571.04 -1.52 571.36 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 572.395 8.675 572.725 9.005 ;
        RECT 572.395 7.315 572.725 7.645 ;
        RECT 572.395 1.875 572.725 2.205 ;
        RECT 572.395 0.515 572.725 0.845 ;
        RECT 572.395 -0.845 572.725 -0.515 ;
        RECT 572.4 -1.52 572.72 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 573.755 8.675 574.085 9.005 ;
        RECT 573.755 7.315 574.085 7.645 ;
        RECT 573.755 1.875 574.085 2.205 ;
        RECT 573.755 0.515 574.085 0.845 ;
        RECT 573.755 -0.845 574.085 -0.515 ;
        RECT 573.76 -1.52 574.08 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 575.115 8.675 575.445 9.005 ;
        RECT 575.115 7.315 575.445 7.645 ;
        RECT 575.115 1.875 575.445 2.205 ;
        RECT 575.115 0.515 575.445 0.845 ;
        RECT 575.115 -0.845 575.445 -0.515 ;
        RECT 575.12 -1.52 575.44 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 576.475 8.675 576.805 9.005 ;
        RECT 576.475 7.315 576.805 7.645 ;
        RECT 576.475 1.875 576.805 2.205 ;
        RECT 576.475 0.515 576.805 0.845 ;
        RECT 576.475 -0.845 576.805 -0.515 ;
        RECT 576.48 -1.52 576.8 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 577.835 8.675 578.165 9.005 ;
        RECT 577.835 7.315 578.165 7.645 ;
        RECT 577.835 1.875 578.165 2.205 ;
        RECT 577.835 0.515 578.165 0.845 ;
        RECT 577.835 -0.845 578.165 -0.515 ;
        RECT 577.84 -1.52 578.16 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 579.195 8.675 579.525 9.005 ;
        RECT 579.195 7.315 579.525 7.645 ;
        RECT 579.195 3.235 579.525 3.565 ;
        RECT 579.195 1.875 579.525 2.205 ;
        RECT 579.195 0.515 579.525 0.845 ;
        RECT 579.195 -0.845 579.525 -0.515 ;
        RECT 579.2 -1.52 579.52 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 580.555 8.675 580.885 9.005 ;
        RECT 580.555 7.315 580.885 7.645 ;
        RECT 580.555 3.235 580.885 3.565 ;
        RECT 580.555 1.875 580.885 2.205 ;
        RECT 580.555 0.515 580.885 0.845 ;
        RECT 580.555 -0.845 580.885 -0.515 ;
        RECT 580.56 -1.52 580.88 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 581.915 8.675 582.245 9.005 ;
        RECT 581.915 7.315 582.245 7.645 ;
        RECT 581.915 3.235 582.245 3.565 ;
        RECT 581.915 1.875 582.245 2.205 ;
        RECT 581.915 0.515 582.245 0.845 ;
        RECT 581.915 -0.845 582.245 -0.515 ;
        RECT 581.92 -1.52 582.24 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 583.275 8.675 583.605 9.005 ;
        RECT 583.275 7.315 583.605 7.645 ;
        RECT 583.275 1.875 583.605 2.205 ;
        RECT 583.275 0.515 583.605 0.845 ;
        RECT 583.275 -0.845 583.605 -0.515 ;
        RECT 583.28 -1.52 583.6 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 584.635 8.675 584.965 9.005 ;
        RECT 584.635 7.315 584.965 7.645 ;
        RECT 584.635 1.875 584.965 2.205 ;
        RECT 584.635 0.515 584.965 0.845 ;
        RECT 584.635 -0.845 584.965 -0.515 ;
        RECT 584.64 -1.52 584.96 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 585.995 8.675 586.325 9.005 ;
        RECT 585.995 7.315 586.325 7.645 ;
        RECT 585.995 1.875 586.325 2.205 ;
        RECT 585.995 0.515 586.325 0.845 ;
        RECT 585.995 -0.845 586.325 -0.515 ;
        RECT 586 -1.52 586.32 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 587.355 8.675 587.685 9.005 ;
        RECT 587.355 7.315 587.685 7.645 ;
        RECT 587.355 1.875 587.685 2.205 ;
        RECT 587.355 0.515 587.685 0.845 ;
        RECT 587.355 -0.845 587.685 -0.515 ;
        RECT 587.36 -1.52 587.68 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 588.715 8.675 589.045 9.005 ;
        RECT 588.715 7.315 589.045 7.645 ;
        RECT 588.715 1.875 589.045 2.205 ;
        RECT 588.715 0.515 589.045 0.845 ;
        RECT 588.715 -0.845 589.045 -0.515 ;
        RECT 588.72 -1.52 589.04 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 590.075 8.675 590.405 9.005 ;
        RECT 590.075 7.315 590.405 7.645 ;
        RECT 590.075 1.875 590.405 2.205 ;
        RECT 590.075 0.515 590.405 0.845 ;
        RECT 590.075 -0.845 590.405 -0.515 ;
        RECT 590.08 -1.52 590.4 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 591.435 8.675 591.765 9.005 ;
        RECT 591.435 7.315 591.765 7.645 ;
        RECT 591.435 3.235 591.765 3.565 ;
        RECT 591.435 1.875 591.765 2.205 ;
        RECT 591.435 0.515 591.765 0.845 ;
        RECT 591.435 -0.845 591.765 -0.515 ;
        RECT 591.44 -1.52 591.76 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 592.795 8.675 593.125 9.005 ;
        RECT 592.795 7.315 593.125 7.645 ;
        RECT 592.795 3.235 593.125 3.565 ;
        RECT 592.795 1.875 593.125 2.205 ;
        RECT 592.795 0.515 593.125 0.845 ;
        RECT 592.795 -0.845 593.125 -0.515 ;
        RECT 592.8 -1.52 593.12 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 594.155 8.675 594.485 9.005 ;
        RECT 594.155 7.315 594.485 7.645 ;
        RECT 594.155 3.235 594.485 3.565 ;
        RECT 594.155 1.875 594.485 2.205 ;
        RECT 594.155 0.515 594.485 0.845 ;
        RECT 594.155 -0.845 594.485 -0.515 ;
        RECT 594.16 -1.52 594.48 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 595.515 8.675 595.845 9.005 ;
        RECT 595.515 7.315 595.845 7.645 ;
        RECT 595.515 1.875 595.845 2.205 ;
        RECT 595.515 0.515 595.845 0.845 ;
        RECT 595.515 -0.845 595.845 -0.515 ;
        RECT 595.52 -1.52 595.84 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 596.875 8.675 597.205 9.005 ;
        RECT 596.875 7.315 597.205 7.645 ;
        RECT 596.875 1.875 597.205 2.205 ;
        RECT 596.875 0.515 597.205 0.845 ;
        RECT 596.875 -0.845 597.205 -0.515 ;
        RECT 596.88 -1.52 597.2 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 598.235 8.675 598.565 9.005 ;
        RECT 598.235 7.315 598.565 7.645 ;
        RECT 598.235 1.875 598.565 2.205 ;
        RECT 598.235 0.515 598.565 0.845 ;
        RECT 598.235 -0.845 598.565 -0.515 ;
        RECT 598.24 -1.52 598.56 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 599.595 8.675 599.925 9.005 ;
        RECT 599.595 7.315 599.925 7.645 ;
        RECT 599.595 1.875 599.925 2.205 ;
        RECT 599.595 0.515 599.925 0.845 ;
        RECT 599.595 -0.845 599.925 -0.515 ;
        RECT 599.6 -1.52 599.92 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 600.955 8.675 601.285 9.005 ;
        RECT 600.955 7.315 601.285 7.645 ;
        RECT 600.955 1.875 601.285 2.205 ;
        RECT 600.955 0.515 601.285 0.845 ;
        RECT 600.955 -0.845 601.285 -0.515 ;
        RECT 600.96 -1.52 601.28 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 602.315 8.675 602.645 9.005 ;
        RECT 602.315 7.315 602.645 7.645 ;
        RECT 602.315 1.875 602.645 2.205 ;
        RECT 602.315 0.515 602.645 0.845 ;
        RECT 602.315 -0.845 602.645 -0.515 ;
        RECT 602.32 -1.52 602.64 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 603.675 8.675 604.005 9.005 ;
        RECT 603.675 7.315 604.005 7.645 ;
        RECT 603.675 3.235 604.005 3.565 ;
        RECT 603.675 1.875 604.005 2.205 ;
        RECT 603.675 0.515 604.005 0.845 ;
        RECT 603.675 -0.845 604.005 -0.515 ;
        RECT 603.68 -1.52 604 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 605.035 8.675 605.365 9.005 ;
        RECT 605.035 7.315 605.365 7.645 ;
        RECT 605.035 3.235 605.365 3.565 ;
        RECT 605.035 1.875 605.365 2.205 ;
        RECT 605.035 0.515 605.365 0.845 ;
        RECT 605.035 -0.845 605.365 -0.515 ;
        RECT 605.04 -1.52 605.36 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 606.395 8.675 606.725 9.005 ;
        RECT 606.395 7.315 606.725 7.645 ;
        RECT 606.395 3.235 606.725 3.565 ;
        RECT 606.395 1.875 606.725 2.205 ;
        RECT 606.395 0.515 606.725 0.845 ;
        RECT 606.395 -0.845 606.725 -0.515 ;
        RECT 606.4 -1.52 606.72 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 607.755 8.675 608.085 9.005 ;
        RECT 607.755 7.315 608.085 7.645 ;
        RECT 607.755 1.875 608.085 2.205 ;
        RECT 607.755 0.515 608.085 0.845 ;
        RECT 607.755 -0.845 608.085 -0.515 ;
        RECT 607.76 -1.52 608.08 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 609.115 8.675 609.445 9.005 ;
        RECT 609.115 7.315 609.445 7.645 ;
        RECT 609.115 1.875 609.445 2.205 ;
        RECT 609.115 0.515 609.445 0.845 ;
        RECT 609.115 -0.845 609.445 -0.515 ;
        RECT 609.12 -1.52 609.44 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 610.475 8.675 610.805 9.005 ;
        RECT 610.475 7.315 610.805 7.645 ;
        RECT 610.475 1.875 610.805 2.205 ;
        RECT 610.475 0.515 610.805 0.845 ;
        RECT 610.475 -0.845 610.805 -0.515 ;
        RECT 610.48 -1.52 610.8 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 611.835 8.675 612.165 9.005 ;
        RECT 611.835 7.315 612.165 7.645 ;
        RECT 611.835 1.875 612.165 2.205 ;
        RECT 611.835 0.515 612.165 0.845 ;
        RECT 611.835 -0.845 612.165 -0.515 ;
        RECT 611.84 -1.52 612.16 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 613.195 8.675 613.525 9.005 ;
        RECT 613.195 7.315 613.525 7.645 ;
        RECT 613.195 1.875 613.525 2.205 ;
        RECT 613.195 0.515 613.525 0.845 ;
        RECT 613.195 -0.845 613.525 -0.515 ;
        RECT 613.2 -1.52 613.52 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 614.555 8.675 614.885 9.005 ;
        RECT 614.555 7.315 614.885 7.645 ;
        RECT 614.555 1.875 614.885 2.205 ;
        RECT 614.555 0.515 614.885 0.845 ;
        RECT 614.555 -0.845 614.885 -0.515 ;
        RECT 614.56 -1.52 614.88 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 615.915 8.675 616.245 9.005 ;
        RECT 615.915 7.315 616.245 7.645 ;
        RECT 615.915 3.235 616.245 3.565 ;
        RECT 615.915 1.875 616.245 2.205 ;
        RECT 615.915 0.515 616.245 0.845 ;
        RECT 615.915 -0.845 616.245 -0.515 ;
        RECT 615.92 -1.52 616.24 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 617.275 8.675 617.605 9.005 ;
        RECT 617.275 7.315 617.605 7.645 ;
        RECT 617.275 3.235 617.605 3.565 ;
        RECT 617.275 1.875 617.605 2.205 ;
        RECT 617.275 0.515 617.605 0.845 ;
        RECT 617.275 -0.845 617.605 -0.515 ;
        RECT 617.28 -1.52 617.6 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 618.635 8.675 618.965 9.005 ;
        RECT 618.635 7.315 618.965 7.645 ;
        RECT 618.635 3.235 618.965 3.565 ;
        RECT 618.635 1.875 618.965 2.205 ;
        RECT 618.635 0.515 618.965 0.845 ;
        RECT 618.635 -0.845 618.965 -0.515 ;
        RECT 618.64 -1.52 618.96 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 619.995 8.675 620.325 9.005 ;
        RECT 619.995 7.315 620.325 7.645 ;
        RECT 619.995 1.875 620.325 2.205 ;
        RECT 619.995 0.515 620.325 0.845 ;
        RECT 619.995 -0.845 620.325 -0.515 ;
        RECT 620 -1.52 620.32 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 621.355 8.675 621.685 9.005 ;
        RECT 621.355 7.315 621.685 7.645 ;
        RECT 621.355 1.875 621.685 2.205 ;
        RECT 621.355 0.515 621.685 0.845 ;
        RECT 621.355 -0.845 621.685 -0.515 ;
        RECT 621.36 -1.52 621.68 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 622.715 8.675 623.045 9.005 ;
        RECT 622.715 7.315 623.045 7.645 ;
        RECT 622.715 1.875 623.045 2.205 ;
        RECT 622.715 0.515 623.045 0.845 ;
        RECT 622.715 -0.845 623.045 -0.515 ;
        RECT 622.72 -1.52 623.04 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 624.075 8.675 624.405 9.005 ;
        RECT 624.075 7.315 624.405 7.645 ;
        RECT 624.075 1.875 624.405 2.205 ;
        RECT 624.075 0.515 624.405 0.845 ;
        RECT 624.075 -0.845 624.405 -0.515 ;
        RECT 624.08 -1.52 624.4 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 625.435 8.675 625.765 9.005 ;
        RECT 625.435 7.315 625.765 7.645 ;
        RECT 625.435 1.875 625.765 2.205 ;
        RECT 625.435 0.515 625.765 0.845 ;
        RECT 625.435 -0.845 625.765 -0.515 ;
        RECT 625.44 -1.52 625.76 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 626.795 8.675 627.125 9.005 ;
        RECT 626.795 7.315 627.125 7.645 ;
        RECT 626.795 1.875 627.125 2.205 ;
        RECT 626.795 0.515 627.125 0.845 ;
        RECT 626.795 -0.845 627.125 -0.515 ;
        RECT 626.8 -1.52 627.12 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 628.155 8.675 628.485 9.005 ;
        RECT 628.155 7.315 628.485 7.645 ;
        RECT 628.155 3.235 628.485 3.565 ;
        RECT 628.155 1.875 628.485 2.205 ;
        RECT 628.155 0.515 628.485 0.845 ;
        RECT 628.155 -0.845 628.485 -0.515 ;
        RECT 628.16 -1.52 628.48 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 629.515 8.675 629.845 9.005 ;
        RECT 629.515 7.315 629.845 7.645 ;
        RECT 629.515 3.235 629.845 3.565 ;
        RECT 629.515 1.875 629.845 2.205 ;
        RECT 629.515 0.515 629.845 0.845 ;
        RECT 629.515 -0.845 629.845 -0.515 ;
        RECT 629.52 -1.52 629.84 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 630.875 8.675 631.205 9.005 ;
        RECT 630.875 7.315 631.205 7.645 ;
        RECT 630.875 1.875 631.205 2.205 ;
        RECT 630.875 0.515 631.205 0.845 ;
        RECT 630.875 -0.845 631.205 -0.515 ;
        RECT 630.88 -1.52 631.2 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 632.235 8.675 632.565 9.005 ;
        RECT 632.235 7.315 632.565 7.645 ;
        RECT 632.235 1.875 632.565 2.205 ;
        RECT 632.235 0.515 632.565 0.845 ;
        RECT 632.235 -0.845 632.565 -0.515 ;
        RECT 632.24 -1.52 632.56 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 633.595 8.675 633.925 9.005 ;
        RECT 633.595 7.315 633.925 7.645 ;
        RECT 633.595 1.875 633.925 2.205 ;
        RECT 633.595 0.515 633.925 0.845 ;
        RECT 633.595 -0.845 633.925 -0.515 ;
        RECT 633.6 -1.52 633.92 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 634.955 8.675 635.285 9.005 ;
        RECT 634.955 7.315 635.285 7.645 ;
        RECT 634.955 1.875 635.285 2.205 ;
        RECT 634.955 0.515 635.285 0.845 ;
        RECT 634.955 -0.845 635.285 -0.515 ;
        RECT 634.96 -1.52 635.28 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 636.315 8.675 636.645 9.005 ;
        RECT 636.315 7.315 636.645 7.645 ;
        RECT 636.315 1.875 636.645 2.205 ;
        RECT 636.315 0.515 636.645 0.845 ;
        RECT 636.315 -0.845 636.645 -0.515 ;
        RECT 636.32 -1.52 636.64 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 637.675 8.675 638.005 9.005 ;
        RECT 637.675 7.315 638.005 7.645 ;
        RECT 637.675 1.875 638.005 2.205 ;
        RECT 637.675 0.515 638.005 0.845 ;
        RECT 637.675 -0.845 638.005 -0.515 ;
        RECT 637.68 -1.52 638 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 639.035 8.675 639.365 9.005 ;
        RECT 639.035 7.315 639.365 7.645 ;
        RECT 639.035 3.235 639.365 3.565 ;
        RECT 639.035 1.875 639.365 2.205 ;
        RECT 639.035 0.515 639.365 0.845 ;
        RECT 639.035 -0.845 639.365 -0.515 ;
        RECT 639.04 -1.52 639.36 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 640.395 8.675 640.725 9.005 ;
        RECT 640.395 7.315 640.725 7.645 ;
        RECT 640.395 3.235 640.725 3.565 ;
        RECT 640.395 1.875 640.725 2.205 ;
        RECT 640.395 0.515 640.725 0.845 ;
        RECT 640.395 -0.845 640.725 -0.515 ;
        RECT 640.4 -1.52 640.72 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 641.755 8.675 642.085 9.005 ;
        RECT 641.755 7.315 642.085 7.645 ;
        RECT 641.755 3.235 642.085 3.565 ;
        RECT 641.755 1.875 642.085 2.205 ;
        RECT 641.755 0.515 642.085 0.845 ;
        RECT 641.755 -0.845 642.085 -0.515 ;
        RECT 641.76 -1.52 642.08 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 643.115 8.675 643.445 9.005 ;
        RECT 643.115 7.315 643.445 7.645 ;
        RECT 643.115 1.875 643.445 2.205 ;
        RECT 643.115 0.515 643.445 0.845 ;
        RECT 643.115 -0.845 643.445 -0.515 ;
        RECT 643.12 -1.52 643.44 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 644.475 8.675 644.805 9.005 ;
        RECT 644.475 7.315 644.805 7.645 ;
        RECT 644.475 1.875 644.805 2.205 ;
        RECT 644.475 0.515 644.805 0.845 ;
        RECT 644.475 -0.845 644.805 -0.515 ;
        RECT 644.48 -1.52 644.8 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 645.835 8.675 646.165 9.005 ;
        RECT 645.835 7.315 646.165 7.645 ;
        RECT 645.835 1.875 646.165 2.205 ;
        RECT 645.835 0.515 646.165 0.845 ;
        RECT 645.835 -0.845 646.165 -0.515 ;
        RECT 645.84 -1.52 646.16 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 647.195 8.675 647.525 9.005 ;
        RECT 647.195 7.315 647.525 7.645 ;
        RECT 647.195 1.875 647.525 2.205 ;
        RECT 647.195 0.515 647.525 0.845 ;
        RECT 647.195 -0.845 647.525 -0.515 ;
        RECT 647.2 -1.52 647.52 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 648.555 8.675 648.885 9.005 ;
        RECT 648.555 7.315 648.885 7.645 ;
        RECT 648.555 1.875 648.885 2.205 ;
        RECT 648.555 0.515 648.885 0.845 ;
        RECT 648.555 -0.845 648.885 -0.515 ;
        RECT 648.56 -1.52 648.88 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 649.915 8.675 650.245 9.005 ;
        RECT 649.915 7.315 650.245 7.645 ;
        RECT 649.915 1.875 650.245 2.205 ;
        RECT 649.915 0.515 650.245 0.845 ;
        RECT 649.915 -0.845 650.245 -0.515 ;
        RECT 649.92 -1.52 650.24 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 651.275 8.675 651.605 9.005 ;
        RECT 651.275 7.315 651.605 7.645 ;
        RECT 651.275 3.235 651.605 3.565 ;
        RECT 651.275 1.875 651.605 2.205 ;
        RECT 651.275 0.515 651.605 0.845 ;
        RECT 651.275 -0.845 651.605 -0.515 ;
        RECT 651.28 -1.52 651.6 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 652.635 8.675 652.965 9.005 ;
        RECT 652.635 7.315 652.965 7.645 ;
        RECT 652.635 3.235 652.965 3.565 ;
        RECT 652.635 1.875 652.965 2.205 ;
        RECT 652.635 0.515 652.965 0.845 ;
        RECT 652.635 -0.845 652.965 -0.515 ;
        RECT 652.64 -1.52 652.96 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 653.995 8.675 654.325 9.005 ;
        RECT 653.995 7.315 654.325 7.645 ;
        RECT 653.995 3.235 654.325 3.565 ;
        RECT 653.995 1.875 654.325 2.205 ;
        RECT 653.995 0.515 654.325 0.845 ;
        RECT 653.995 -0.845 654.325 -0.515 ;
        RECT 654 -1.52 654.32 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 655.355 8.675 655.685 9.005 ;
        RECT 655.355 7.315 655.685 7.645 ;
        RECT 655.355 1.875 655.685 2.205 ;
        RECT 655.355 0.515 655.685 0.845 ;
        RECT 655.355 -0.845 655.685 -0.515 ;
        RECT 655.36 -1.52 655.68 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 656.715 8.675 657.045 9.005 ;
        RECT 656.715 7.315 657.045 7.645 ;
        RECT 656.715 1.875 657.045 2.205 ;
        RECT 656.715 0.515 657.045 0.845 ;
        RECT 656.715 -0.845 657.045 -0.515 ;
        RECT 656.72 -1.52 657.04 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 658.075 8.675 658.405 9.005 ;
        RECT 658.075 7.315 658.405 7.645 ;
        RECT 658.075 1.875 658.405 2.205 ;
        RECT 658.075 0.515 658.405 0.845 ;
        RECT 658.075 -0.845 658.405 -0.515 ;
        RECT 658.08 -1.52 658.4 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 659.435 8.675 659.765 9.005 ;
        RECT 659.435 7.315 659.765 7.645 ;
        RECT 659.435 1.875 659.765 2.205 ;
        RECT 659.435 0.515 659.765 0.845 ;
        RECT 659.435 -0.845 659.765 -0.515 ;
        RECT 659.44 -1.52 659.76 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 660.795 8.675 661.125 9.005 ;
        RECT 660.795 7.315 661.125 7.645 ;
        RECT 660.795 1.875 661.125 2.205 ;
        RECT 660.795 0.515 661.125 0.845 ;
        RECT 660.795 -0.845 661.125 -0.515 ;
        RECT 660.8 -1.52 661.12 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 662.155 8.675 662.485 9.005 ;
        RECT 662.155 7.315 662.485 7.645 ;
        RECT 662.155 1.875 662.485 2.205 ;
        RECT 662.155 0.515 662.485 0.845 ;
        RECT 662.155 -0.845 662.485 -0.515 ;
        RECT 662.16 -1.52 662.48 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 663.515 8.675 663.845 9.005 ;
        RECT 663.515 7.315 663.845 7.645 ;
        RECT 663.515 3.235 663.845 3.565 ;
        RECT 663.515 1.875 663.845 2.205 ;
        RECT 663.515 0.515 663.845 0.845 ;
        RECT 663.515 -0.845 663.845 -0.515 ;
        RECT 663.52 -1.52 663.84 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 664.875 8.675 665.205 9.005 ;
        RECT 664.875 7.315 665.205 7.645 ;
        RECT 664.875 3.235 665.205 3.565 ;
        RECT 664.875 1.875 665.205 2.205 ;
        RECT 664.875 0.515 665.205 0.845 ;
        RECT 664.875 -0.845 665.205 -0.515 ;
        RECT 664.88 -1.52 665.2 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 666.235 8.675 666.565 9.005 ;
        RECT 666.235 7.315 666.565 7.645 ;
        RECT 666.235 3.235 666.565 3.565 ;
        RECT 666.235 1.875 666.565 2.205 ;
        RECT 666.235 0.515 666.565 0.845 ;
        RECT 666.235 -0.845 666.565 -0.515 ;
        RECT 666.24 -1.52 666.56 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 667.595 8.675 667.925 9.005 ;
        RECT 667.595 7.315 667.925 7.645 ;
        RECT 667.595 1.875 667.925 2.205 ;
        RECT 667.595 0.515 667.925 0.845 ;
        RECT 667.595 -0.845 667.925 -0.515 ;
        RECT 667.6 -1.52 667.92 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 668.955 8.675 669.285 9.005 ;
        RECT 668.955 7.315 669.285 7.645 ;
        RECT 668.955 1.875 669.285 2.205 ;
        RECT 668.955 0.515 669.285 0.845 ;
        RECT 668.955 -0.845 669.285 -0.515 ;
        RECT 668.96 -1.52 669.28 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 670.315 8.675 670.645 9.005 ;
        RECT 670.315 7.315 670.645 7.645 ;
        RECT 670.315 1.875 670.645 2.205 ;
        RECT 670.315 0.515 670.645 0.845 ;
        RECT 670.315 -0.845 670.645 -0.515 ;
        RECT 670.32 -1.52 670.64 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 671.675 8.675 672.005 9.005 ;
        RECT 671.675 7.315 672.005 7.645 ;
        RECT 671.675 1.875 672.005 2.205 ;
        RECT 671.675 0.515 672.005 0.845 ;
        RECT 671.675 -0.845 672.005 -0.515 ;
        RECT 671.68 -1.52 672 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 673.035 8.675 673.365 9.005 ;
        RECT 673.035 7.315 673.365 7.645 ;
        RECT 673.035 1.875 673.365 2.205 ;
        RECT 673.035 0.515 673.365 0.845 ;
        RECT 673.035 -0.845 673.365 -0.515 ;
        RECT 673.04 -1.52 673.36 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 674.395 8.675 674.725 9.005 ;
        RECT 674.395 7.315 674.725 7.645 ;
        RECT 674.395 1.875 674.725 2.205 ;
        RECT 674.395 0.515 674.725 0.845 ;
        RECT 674.395 -0.845 674.725 -0.515 ;
        RECT 674.4 -1.52 674.72 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 675.755 8.675 676.085 9.005 ;
        RECT 675.755 7.315 676.085 7.645 ;
        RECT 675.755 3.235 676.085 3.565 ;
        RECT 675.755 1.875 676.085 2.205 ;
        RECT 675.755 0.515 676.085 0.845 ;
        RECT 675.755 -0.845 676.085 -0.515 ;
        RECT 675.76 -1.52 676.08 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 677.115 8.675 677.445 9.005 ;
        RECT 677.115 7.315 677.445 7.645 ;
        RECT 677.115 3.235 677.445 3.565 ;
        RECT 677.115 1.875 677.445 2.205 ;
        RECT 677.115 0.515 677.445 0.845 ;
        RECT 677.115 -0.845 677.445 -0.515 ;
        RECT 677.12 -1.52 677.44 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 678.475 8.675 678.805 9.005 ;
        RECT 678.475 7.315 678.805 7.645 ;
        RECT 678.475 3.235 678.805 3.565 ;
        RECT 678.475 1.875 678.805 2.205 ;
        RECT 678.475 0.515 678.805 0.845 ;
        RECT 678.475 -0.845 678.805 -0.515 ;
        RECT 678.48 -1.52 678.8 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 679.835 8.675 680.165 9.005 ;
        RECT 679.835 7.315 680.165 7.645 ;
        RECT 679.835 1.875 680.165 2.205 ;
        RECT 679.835 0.515 680.165 0.845 ;
        RECT 679.835 -0.845 680.165 -0.515 ;
        RECT 679.84 -1.52 680.16 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 681.195 8.675 681.525 9.005 ;
        RECT 681.195 7.315 681.525 7.645 ;
        RECT 681.195 1.875 681.525 2.205 ;
        RECT 681.195 0.515 681.525 0.845 ;
        RECT 681.195 -0.845 681.525 -0.515 ;
        RECT 681.2 -1.52 681.52 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 682.555 8.675 682.885 9.005 ;
        RECT 682.555 7.315 682.885 7.645 ;
        RECT 682.555 1.875 682.885 2.205 ;
        RECT 682.555 0.515 682.885 0.845 ;
        RECT 682.555 -0.845 682.885 -0.515 ;
        RECT 682.56 -1.52 682.88 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 683.915 8.675 684.245 9.005 ;
        RECT 683.915 7.315 684.245 7.645 ;
        RECT 683.915 1.875 684.245 2.205 ;
        RECT 683.915 0.515 684.245 0.845 ;
        RECT 683.915 -0.845 684.245 -0.515 ;
        RECT 683.92 -1.52 684.24 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 685.275 8.675 685.605 9.005 ;
        RECT 685.275 7.315 685.605 7.645 ;
        RECT 685.275 1.875 685.605 2.205 ;
        RECT 685.275 0.515 685.605 0.845 ;
        RECT 685.275 -0.845 685.605 -0.515 ;
        RECT 685.28 -1.52 685.6 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 686.635 8.675 686.965 9.005 ;
        RECT 686.635 7.315 686.965 7.645 ;
        RECT 686.635 1.875 686.965 2.205 ;
        RECT 686.635 0.515 686.965 0.845 ;
        RECT 686.635 -0.845 686.965 -0.515 ;
        RECT 686.64 -1.52 686.96 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 687.995 8.675 688.325 9.005 ;
        RECT 687.995 7.315 688.325 7.645 ;
        RECT 687.995 3.235 688.325 3.565 ;
        RECT 687.995 1.875 688.325 2.205 ;
        RECT 687.995 0.515 688.325 0.845 ;
        RECT 687.995 -0.845 688.325 -0.515 ;
        RECT 688 -1.52 688.32 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 689.355 8.675 689.685 9.005 ;
        RECT 689.355 7.315 689.685 7.645 ;
        RECT 689.355 3.235 689.685 3.565 ;
        RECT 689.355 1.875 689.685 2.205 ;
        RECT 689.355 0.515 689.685 0.845 ;
        RECT 689.355 -0.845 689.685 -0.515 ;
        RECT 689.36 -1.52 689.68 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 690.715 8.675 691.045 9.005 ;
        RECT 690.715 7.315 691.045 7.645 ;
        RECT 690.715 3.235 691.045 3.565 ;
        RECT 690.715 1.875 691.045 2.205 ;
        RECT 690.715 0.515 691.045 0.845 ;
        RECT 690.715 -0.845 691.045 -0.515 ;
        RECT 690.72 -1.52 691.04 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 692.075 8.675 692.405 9.005 ;
        RECT 692.075 7.315 692.405 7.645 ;
        RECT 692.075 1.875 692.405 2.205 ;
        RECT 692.075 0.515 692.405 0.845 ;
        RECT 692.075 -0.845 692.405 -0.515 ;
        RECT 692.08 -1.52 692.4 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 693.435 8.675 693.765 9.005 ;
        RECT 693.435 7.315 693.765 7.645 ;
        RECT 693.435 1.875 693.765 2.205 ;
        RECT 693.435 0.515 693.765 0.845 ;
        RECT 693.435 -0.845 693.765 -0.515 ;
        RECT 693.44 -1.52 693.76 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 694.795 8.675 695.125 9.005 ;
        RECT 694.795 7.315 695.125 7.645 ;
        RECT 694.795 1.875 695.125 2.205 ;
        RECT 694.795 0.515 695.125 0.845 ;
        RECT 694.795 -0.845 695.125 -0.515 ;
        RECT 694.8 -1.52 695.12 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 696.155 8.675 696.485 9.005 ;
        RECT 696.155 7.315 696.485 7.645 ;
        RECT 696.155 1.875 696.485 2.205 ;
        RECT 696.155 0.515 696.485 0.845 ;
        RECT 696.155 -0.845 696.485 -0.515 ;
        RECT 696.16 -1.52 696.48 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 697.515 8.675 697.845 9.005 ;
        RECT 697.515 7.315 697.845 7.645 ;
        RECT 697.515 1.875 697.845 2.205 ;
        RECT 697.515 0.515 697.845 0.845 ;
        RECT 697.515 -0.845 697.845 -0.515 ;
        RECT 697.52 -1.52 697.84 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 698.875 8.675 699.205 9.005 ;
        RECT 698.875 7.315 699.205 7.645 ;
        RECT 698.875 3.235 699.205 3.565 ;
        RECT 698.875 1.875 699.205 2.205 ;
        RECT 698.875 0.515 699.205 0.845 ;
        RECT 698.875 -0.845 699.205 -0.515 ;
        RECT 698.88 -1.52 699.2 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 700.235 8.675 700.565 9.005 ;
        RECT 700.235 7.315 700.565 7.645 ;
        RECT 700.235 3.235 700.565 3.565 ;
        RECT 700.235 1.875 700.565 2.205 ;
        RECT 700.235 0.515 700.565 0.845 ;
        RECT 700.235 -0.845 700.565 -0.515 ;
        RECT 700.24 -1.52 700.56 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 701.595 8.675 701.925 9.005 ;
        RECT 701.595 7.315 701.925 7.645 ;
        RECT 701.595 3.235 701.925 3.565 ;
        RECT 701.595 1.875 701.925 2.205 ;
        RECT 701.595 0.515 701.925 0.845 ;
        RECT 701.595 -0.845 701.925 -0.515 ;
        RECT 701.6 -1.52 701.92 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 702.955 8.675 703.285 9.005 ;
        RECT 702.955 7.315 703.285 7.645 ;
        RECT 702.955 1.875 703.285 2.205 ;
        RECT 702.955 0.515 703.285 0.845 ;
        RECT 702.955 -0.845 703.285 -0.515 ;
        RECT 702.96 -1.52 703.28 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 704.315 8.675 704.645 9.005 ;
        RECT 704.315 7.315 704.645 7.645 ;
        RECT 704.315 1.875 704.645 2.205 ;
        RECT 704.315 0.515 704.645 0.845 ;
        RECT 704.315 -0.845 704.645 -0.515 ;
        RECT 704.32 -1.52 704.64 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 705.675 8.675 706.005 9.005 ;
        RECT 705.675 7.315 706.005 7.645 ;
        RECT 705.675 1.875 706.005 2.205 ;
        RECT 705.675 0.515 706.005 0.845 ;
        RECT 705.675 -0.845 706.005 -0.515 ;
        RECT 705.68 -1.52 706 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 707.035 8.675 707.365 9.005 ;
        RECT 707.035 7.315 707.365 7.645 ;
        RECT 707.035 1.875 707.365 2.205 ;
        RECT 707.035 0.515 707.365 0.845 ;
        RECT 707.035 -0.845 707.365 -0.515 ;
        RECT 707.04 -1.52 707.36 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 708.395 8.675 708.725 9.005 ;
        RECT 708.395 7.315 708.725 7.645 ;
        RECT 708.395 1.875 708.725 2.205 ;
        RECT 708.395 0.515 708.725 0.845 ;
        RECT 708.395 -0.845 708.725 -0.515 ;
        RECT 708.4 -1.52 708.72 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 709.755 8.675 710.085 9.005 ;
        RECT 709.755 7.315 710.085 7.645 ;
        RECT 709.755 1.875 710.085 2.205 ;
        RECT 709.755 0.515 710.085 0.845 ;
        RECT 709.755 -0.845 710.085 -0.515 ;
        RECT 709.76 -1.52 710.08 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 711.115 8.675 711.445 9.005 ;
        RECT 711.115 7.315 711.445 7.645 ;
        RECT 711.115 3.235 711.445 3.565 ;
        RECT 711.115 1.875 711.445 2.205 ;
        RECT 711.115 0.515 711.445 0.845 ;
        RECT 711.115 -0.845 711.445 -0.515 ;
        RECT 711.12 -1.52 711.44 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 712.475 8.675 712.805 9.005 ;
        RECT 712.475 7.315 712.805 7.645 ;
        RECT 712.475 3.235 712.805 3.565 ;
        RECT 712.475 1.875 712.805 2.205 ;
        RECT 712.475 0.515 712.805 0.845 ;
        RECT 712.475 -0.845 712.805 -0.515 ;
        RECT 712.48 -1.52 712.8 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 713.835 8.675 714.165 9.005 ;
        RECT 713.835 7.315 714.165 7.645 ;
        RECT 713.835 3.235 714.165 3.565 ;
        RECT 713.835 1.875 714.165 2.205 ;
        RECT 713.835 0.515 714.165 0.845 ;
        RECT 713.835 -0.845 714.165 -0.515 ;
        RECT 713.84 -1.52 714.16 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 715.195 8.675 715.525 9.005 ;
        RECT 715.195 7.315 715.525 7.645 ;
        RECT 715.195 1.875 715.525 2.205 ;
        RECT 715.195 0.515 715.525 0.845 ;
        RECT 715.195 -0.845 715.525 -0.515 ;
        RECT 715.2 -1.52 715.52 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 716.555 8.675 716.885 9.005 ;
        RECT 716.555 7.315 716.885 7.645 ;
        RECT 716.555 1.875 716.885 2.205 ;
        RECT 716.555 0.515 716.885 0.845 ;
        RECT 716.555 -0.845 716.885 -0.515 ;
        RECT 716.56 -1.52 716.88 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 717.915 8.675 718.245 9.005 ;
        RECT 717.915 7.315 718.245 7.645 ;
        RECT 717.915 1.875 718.245 2.205 ;
        RECT 717.915 0.515 718.245 0.845 ;
        RECT 717.915 -0.845 718.245 -0.515 ;
        RECT 717.92 -1.52 718.24 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 719.275 8.675 719.605 9.005 ;
        RECT 719.275 7.315 719.605 7.645 ;
        RECT 719.275 1.875 719.605 2.205 ;
        RECT 719.275 0.515 719.605 0.845 ;
        RECT 719.275 -0.845 719.605 -0.515 ;
        RECT 719.28 -1.52 719.6 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 720.635 8.675 720.965 9.005 ;
        RECT 720.635 7.315 720.965 7.645 ;
        RECT 720.635 1.875 720.965 2.205 ;
        RECT 720.635 0.515 720.965 0.845 ;
        RECT 720.635 -0.845 720.965 -0.515 ;
        RECT 720.64 -1.52 720.96 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 721.995 8.675 722.325 9.005 ;
        RECT 721.995 7.315 722.325 7.645 ;
        RECT 721.995 1.875 722.325 2.205 ;
        RECT 721.995 0.515 722.325 0.845 ;
        RECT 721.995 -0.845 722.325 -0.515 ;
        RECT 722 -1.52 722.32 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 723.355 8.675 723.685 9.005 ;
        RECT 723.355 7.315 723.685 7.645 ;
        RECT 723.355 3.235 723.685 3.565 ;
        RECT 723.355 1.875 723.685 2.205 ;
        RECT 723.355 0.515 723.685 0.845 ;
        RECT 723.355 -0.845 723.685 -0.515 ;
        RECT 723.36 -1.52 723.68 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 724.715 8.675 725.045 9.005 ;
        RECT 724.715 7.315 725.045 7.645 ;
        RECT 724.715 3.235 725.045 3.565 ;
        RECT 724.715 1.875 725.045 2.205 ;
        RECT 724.715 0.515 725.045 0.845 ;
        RECT 724.715 -0.845 725.045 -0.515 ;
        RECT 724.72 -1.52 725.04 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 726.075 8.675 726.405 9.005 ;
        RECT 726.075 7.315 726.405 7.645 ;
        RECT 726.075 3.235 726.405 3.565 ;
        RECT 726.075 1.875 726.405 2.205 ;
        RECT 726.075 0.515 726.405 0.845 ;
        RECT 726.075 -0.845 726.405 -0.515 ;
        RECT 726.08 -1.52 726.4 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 727.435 8.675 727.765 9.005 ;
        RECT 727.435 7.315 727.765 7.645 ;
        RECT 727.435 1.875 727.765 2.205 ;
        RECT 727.435 0.515 727.765 0.845 ;
        RECT 727.435 -0.845 727.765 -0.515 ;
        RECT 727.44 -1.52 727.76 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 728.795 8.675 729.125 9.005 ;
        RECT 728.795 7.315 729.125 7.645 ;
        RECT 728.795 1.875 729.125 2.205 ;
        RECT 728.795 0.515 729.125 0.845 ;
        RECT 728.795 -0.845 729.125 -0.515 ;
        RECT 728.8 -1.52 729.12 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 730.155 8.675 730.485 9.005 ;
        RECT 730.155 7.315 730.485 7.645 ;
        RECT 730.155 1.875 730.485 2.205 ;
        RECT 730.155 0.515 730.485 0.845 ;
        RECT 730.155 -0.845 730.485 -0.515 ;
        RECT 730.16 -1.52 730.48 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 731.515 8.675 731.845 9.005 ;
        RECT 731.515 7.315 731.845 7.645 ;
        RECT 731.515 1.875 731.845 2.205 ;
        RECT 731.515 0.515 731.845 0.845 ;
        RECT 731.515 -0.845 731.845 -0.515 ;
        RECT 731.52 -1.52 731.84 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 732.875 8.675 733.205 9.005 ;
        RECT 732.875 7.315 733.205 7.645 ;
        RECT 732.875 1.875 733.205 2.205 ;
        RECT 732.875 0.515 733.205 0.845 ;
        RECT 732.875 -0.845 733.205 -0.515 ;
        RECT 732.88 -1.52 733.2 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 734.235 8.675 734.565 9.005 ;
        RECT 734.235 7.315 734.565 7.645 ;
        RECT 734.235 1.875 734.565 2.205 ;
        RECT 734.235 0.515 734.565 0.845 ;
        RECT 734.235 -0.845 734.565 -0.515 ;
        RECT 734.24 -1.52 734.56 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 735.595 8.675 735.925 9.005 ;
        RECT 735.595 7.315 735.925 7.645 ;
        RECT 735.595 3.235 735.925 3.565 ;
        RECT 735.595 1.875 735.925 2.205 ;
        RECT 735.595 0.515 735.925 0.845 ;
        RECT 735.595 -0.845 735.925 -0.515 ;
        RECT 735.6 -1.52 735.92 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 736.955 8.675 737.285 9.005 ;
        RECT 736.955 7.315 737.285 7.645 ;
        RECT 736.955 3.235 737.285 3.565 ;
        RECT 736.955 1.875 737.285 2.205 ;
        RECT 736.955 0.515 737.285 0.845 ;
        RECT 736.955 -0.845 737.285 -0.515 ;
        RECT 736.96 -1.52 737.28 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 738.315 8.675 738.645 9.005 ;
        RECT 738.315 7.315 738.645 7.645 ;
        RECT 738.315 3.235 738.645 3.565 ;
        RECT 738.315 1.875 738.645 2.205 ;
        RECT 738.315 0.515 738.645 0.845 ;
        RECT 738.315 -0.845 738.645 -0.515 ;
        RECT 738.32 -1.52 738.64 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 739.675 8.675 740.005 9.005 ;
        RECT 739.675 7.315 740.005 7.645 ;
        RECT 739.675 1.875 740.005 2.205 ;
        RECT 739.675 0.515 740.005 0.845 ;
        RECT 739.675 -0.845 740.005 -0.515 ;
        RECT 739.68 -1.52 740 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 741.035 8.675 741.365 9.005 ;
        RECT 741.035 7.315 741.365 7.645 ;
        RECT 741.035 1.875 741.365 2.205 ;
        RECT 741.035 0.515 741.365 0.845 ;
        RECT 741.035 -0.845 741.365 -0.515 ;
        RECT 741.04 -1.52 741.36 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 742.395 8.675 742.725 9.005 ;
        RECT 742.395 7.315 742.725 7.645 ;
        RECT 742.395 1.875 742.725 2.205 ;
        RECT 742.395 0.515 742.725 0.845 ;
        RECT 742.395 -0.845 742.725 -0.515 ;
        RECT 742.4 -1.52 742.72 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 743.755 8.675 744.085 9.005 ;
        RECT 743.755 7.315 744.085 7.645 ;
        RECT 743.755 1.875 744.085 2.205 ;
        RECT 743.755 0.515 744.085 0.845 ;
        RECT 743.755 -0.845 744.085 -0.515 ;
        RECT 743.76 -1.52 744.08 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 745.115 8.675 745.445 9.005 ;
        RECT 745.115 7.315 745.445 7.645 ;
        RECT 745.115 1.875 745.445 2.205 ;
        RECT 745.115 0.515 745.445 0.845 ;
        RECT 745.115 -0.845 745.445 -0.515 ;
        RECT 745.12 -1.52 745.44 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 746.475 8.675 746.805 9.005 ;
        RECT 746.475 7.315 746.805 7.645 ;
        RECT 746.475 1.875 746.805 2.205 ;
        RECT 746.475 0.515 746.805 0.845 ;
        RECT 746.475 -0.845 746.805 -0.515 ;
        RECT 746.48 -1.52 746.8 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 747.835 8.675 748.165 9.005 ;
        RECT 747.835 7.315 748.165 7.645 ;
        RECT 747.835 3.235 748.165 3.565 ;
        RECT 747.835 1.875 748.165 2.205 ;
        RECT 747.835 0.515 748.165 0.845 ;
        RECT 747.835 -0.845 748.165 -0.515 ;
        RECT 747.84 -1.52 748.16 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 749.195 8.675 749.525 9.005 ;
        RECT 749.195 7.315 749.525 7.645 ;
        RECT 749.195 3.235 749.525 3.565 ;
        RECT 749.195 1.875 749.525 2.205 ;
        RECT 749.195 0.515 749.525 0.845 ;
        RECT 749.195 -0.845 749.525 -0.515 ;
        RECT 749.2 -1.52 749.52 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 750.555 8.675 750.885 9.005 ;
        RECT 750.555 7.315 750.885 7.645 ;
        RECT 750.555 3.235 750.885 3.565 ;
        RECT 750.555 1.875 750.885 2.205 ;
        RECT 750.555 0.515 750.885 0.845 ;
        RECT 750.555 -0.845 750.885 -0.515 ;
        RECT 750.56 -1.52 750.88 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 751.915 8.675 752.245 9.005 ;
        RECT 751.915 7.315 752.245 7.645 ;
        RECT 751.915 1.875 752.245 2.205 ;
        RECT 751.915 0.515 752.245 0.845 ;
        RECT 751.915 -0.845 752.245 -0.515 ;
        RECT 751.92 -1.52 752.24 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 753.275 8.675 753.605 9.005 ;
        RECT 753.275 7.315 753.605 7.645 ;
        RECT 753.275 1.875 753.605 2.205 ;
        RECT 753.275 0.515 753.605 0.845 ;
        RECT 753.275 -0.845 753.605 -0.515 ;
        RECT 753.28 -1.52 753.6 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 754.635 8.675 754.965 9.005 ;
        RECT 754.635 7.315 754.965 7.645 ;
        RECT 754.635 1.875 754.965 2.205 ;
        RECT 754.635 0.515 754.965 0.845 ;
        RECT 754.635 -0.845 754.965 -0.515 ;
        RECT 754.64 -1.52 754.96 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 755.995 8.675 756.325 9.005 ;
        RECT 755.995 7.315 756.325 7.645 ;
        RECT 755.995 1.875 756.325 2.205 ;
        RECT 755.995 0.515 756.325 0.845 ;
        RECT 755.995 -0.845 756.325 -0.515 ;
        RECT 756 -1.52 756.32 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 757.355 8.675 757.685 9.005 ;
        RECT 757.355 7.315 757.685 7.645 ;
        RECT 757.355 1.875 757.685 2.205 ;
        RECT 757.355 0.515 757.685 0.845 ;
        RECT 757.355 -0.845 757.685 -0.515 ;
        RECT 757.36 -1.52 757.68 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 758.715 8.675 759.045 9.005 ;
        RECT 758.715 7.315 759.045 7.645 ;
        RECT 758.715 1.875 759.045 2.205 ;
        RECT 758.715 0.515 759.045 0.845 ;
        RECT 758.715 -0.845 759.045 -0.515 ;
        RECT 758.72 -1.52 759.04 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 760.075 8.675 760.405 9.005 ;
        RECT 760.075 7.315 760.405 7.645 ;
        RECT 760.075 3.235 760.405 3.565 ;
        RECT 760.075 1.875 760.405 2.205 ;
        RECT 760.075 0.515 760.405 0.845 ;
        RECT 760.075 -0.845 760.405 -0.515 ;
        RECT 760.08 -1.52 760.4 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 761.435 8.675 761.765 9.005 ;
        RECT 761.435 7.315 761.765 7.645 ;
        RECT 761.435 3.235 761.765 3.565 ;
        RECT 761.435 1.875 761.765 2.205 ;
        RECT 761.435 0.515 761.765 0.845 ;
        RECT 761.435 -0.845 761.765 -0.515 ;
        RECT 761.44 -1.52 761.76 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 762.795 8.675 763.125 9.005 ;
        RECT 762.795 7.315 763.125 7.645 ;
        RECT 762.795 3.235 763.125 3.565 ;
        RECT 762.795 1.875 763.125 2.205 ;
        RECT 762.795 0.515 763.125 0.845 ;
        RECT 762.795 -0.845 763.125 -0.515 ;
        RECT 762.8 -1.52 763.12 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 764.155 8.675 764.485 9.005 ;
        RECT 764.155 7.315 764.485 7.645 ;
        RECT 764.155 3.235 764.485 3.565 ;
        RECT 764.155 1.875 764.485 2.205 ;
        RECT 764.155 0.515 764.485 0.845 ;
        RECT 764.155 -0.845 764.485 -0.515 ;
        RECT 764.16 -1.52 764.48 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 765.515 8.675 765.845 9.005 ;
        RECT 765.515 7.315 765.845 7.645 ;
        RECT 765.515 4.595 765.845 4.925 ;
        RECT 765.515 3.235 765.845 3.565 ;
        RECT 765.515 1.875 765.845 2.205 ;
        RECT 765.515 0.515 765.845 0.845 ;
        RECT 765.515 -0.845 765.845 -0.515 ;
        RECT 765.52 -1.52 765.84 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 766.875 8.675 767.205 9.005 ;
        RECT 766.875 7.315 767.205 7.645 ;
        RECT 766.875 4.595 767.205 4.925 ;
        RECT 766.875 3.235 767.205 3.565 ;
        RECT 766.875 1.875 767.205 2.205 ;
        RECT 766.875 0.515 767.205 0.845 ;
        RECT 766.875 -0.845 767.205 -0.515 ;
        RECT 766.88 -1.52 767.2 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 768.235 8.675 768.565 9.005 ;
        RECT 768.235 7.315 768.565 7.645 ;
        RECT 768.235 5.955 768.565 6.285 ;
        RECT 768.235 4.595 768.565 4.925 ;
        RECT 768.235 3.235 768.565 3.565 ;
        RECT 768.235 1.875 768.565 2.205 ;
        RECT 768.235 0.515 768.565 0.845 ;
        RECT 768.235 -0.845 768.565 -0.515 ;
        RECT 768.24 -1.52 768.56 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 342.555 8.675 342.885 9.005 ;
        RECT 342.555 7.315 342.885 7.645 ;
        RECT 342.555 3.235 342.885 3.565 ;
        RECT 342.555 1.875 342.885 2.205 ;
        RECT 342.555 0.515 342.885 0.845 ;
        RECT 342.555 -0.845 342.885 -0.515 ;
        RECT 342.56 -1.52 342.88 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 343.915 8.675 344.245 9.005 ;
        RECT 343.915 7.315 344.245 7.645 ;
        RECT 343.915 1.875 344.245 2.205 ;
        RECT 343.915 0.515 344.245 0.845 ;
        RECT 343.915 -0.845 344.245 -0.515 ;
        RECT 343.92 -1.52 344.24 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 345.275 8.675 345.605 9.005 ;
        RECT 345.275 7.315 345.605 7.645 ;
        RECT 345.275 1.875 345.605 2.205 ;
        RECT 345.275 0.515 345.605 0.845 ;
        RECT 345.275 -0.845 345.605 -0.515 ;
        RECT 345.28 -1.52 345.6 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 346.635 8.675 346.965 9.005 ;
        RECT 346.635 7.315 346.965 7.645 ;
        RECT 346.635 1.875 346.965 2.205 ;
        RECT 346.635 0.515 346.965 0.845 ;
        RECT 346.635 -0.845 346.965 -0.515 ;
        RECT 346.64 -1.52 346.96 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 347.995 8.675 348.325 9.005 ;
        RECT 347.995 7.315 348.325 7.645 ;
        RECT 347.995 1.875 348.325 2.205 ;
        RECT 347.995 0.515 348.325 0.845 ;
        RECT 347.995 -0.845 348.325 -0.515 ;
        RECT 348 -1.52 348.32 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 349.355 8.675 349.685 9.005 ;
        RECT 349.355 7.315 349.685 7.645 ;
        RECT 349.355 1.875 349.685 2.205 ;
        RECT 349.355 0.515 349.685 0.845 ;
        RECT 349.355 -0.845 349.685 -0.515 ;
        RECT 349.36 -1.52 349.68 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 350.715 8.675 351.045 9.005 ;
        RECT 350.715 7.315 351.045 7.645 ;
        RECT 350.715 1.875 351.045 2.205 ;
        RECT 350.715 0.515 351.045 0.845 ;
        RECT 350.715 -0.845 351.045 -0.515 ;
        RECT 350.72 -1.52 351.04 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 352.075 8.675 352.405 9.005 ;
        RECT 352.075 7.315 352.405 7.645 ;
        RECT 352.075 3.235 352.405 3.565 ;
        RECT 352.075 1.875 352.405 2.205 ;
        RECT 352.075 0.515 352.405 0.845 ;
        RECT 352.075 -0.845 352.405 -0.515 ;
        RECT 352.08 -1.52 352.4 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 353.435 8.675 353.765 9.005 ;
        RECT 353.435 7.315 353.765 7.645 ;
        RECT 353.435 3.235 353.765 3.565 ;
        RECT 353.435 1.875 353.765 2.205 ;
        RECT 353.435 0.515 353.765 0.845 ;
        RECT 353.435 -0.845 353.765 -0.515 ;
        RECT 353.44 -1.52 353.76 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.795 8.675 355.125 9.005 ;
        RECT 354.795 7.315 355.125 7.645 ;
        RECT 354.795 3.235 355.125 3.565 ;
        RECT 354.795 1.875 355.125 2.205 ;
        RECT 354.795 0.515 355.125 0.845 ;
        RECT 354.795 -0.845 355.125 -0.515 ;
        RECT 354.8 -1.52 355.12 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 356.155 8.675 356.485 9.005 ;
        RECT 356.155 7.315 356.485 7.645 ;
        RECT 356.155 1.875 356.485 2.205 ;
        RECT 356.155 0.515 356.485 0.845 ;
        RECT 356.155 -0.845 356.485 -0.515 ;
        RECT 356.16 -1.52 356.48 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 357.515 8.675 357.845 9.005 ;
        RECT 357.515 7.315 357.845 7.645 ;
        RECT 357.515 1.875 357.845 2.205 ;
        RECT 357.515 0.515 357.845 0.845 ;
        RECT 357.515 -0.845 357.845 -0.515 ;
        RECT 357.52 -1.52 357.84 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 358.875 8.675 359.205 9.005 ;
        RECT 358.875 7.315 359.205 7.645 ;
        RECT 358.875 1.875 359.205 2.205 ;
        RECT 358.875 0.515 359.205 0.845 ;
        RECT 358.875 -0.845 359.205 -0.515 ;
        RECT 358.88 -1.52 359.2 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 360.235 8.675 360.565 9.005 ;
        RECT 360.235 7.315 360.565 7.645 ;
        RECT 360.235 1.875 360.565 2.205 ;
        RECT 360.235 0.515 360.565 0.845 ;
        RECT 360.235 -0.845 360.565 -0.515 ;
        RECT 360.24 -1.52 360.56 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 361.595 8.675 361.925 9.005 ;
        RECT 361.595 7.315 361.925 7.645 ;
        RECT 361.595 1.875 361.925 2.205 ;
        RECT 361.595 0.515 361.925 0.845 ;
        RECT 361.595 -0.845 361.925 -0.515 ;
        RECT 361.6 -1.52 361.92 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 362.955 8.675 363.285 9.005 ;
        RECT 362.955 7.315 363.285 7.645 ;
        RECT 362.955 3.235 363.285 3.565 ;
        RECT 362.955 1.875 363.285 2.205 ;
        RECT 362.955 0.515 363.285 0.845 ;
        RECT 362.955 -0.845 363.285 -0.515 ;
        RECT 362.96 -1.52 363.28 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 364.315 8.675 364.645 9.005 ;
        RECT 364.315 7.315 364.645 7.645 ;
        RECT 364.315 3.235 364.645 3.565 ;
        RECT 364.315 1.875 364.645 2.205 ;
        RECT 364.315 0.515 364.645 0.845 ;
        RECT 364.315 -0.845 364.645 -0.515 ;
        RECT 364.32 -1.52 364.64 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 365.675 8.675 366.005 9.005 ;
        RECT 365.675 7.315 366.005 7.645 ;
        RECT 365.675 3.235 366.005 3.565 ;
        RECT 365.675 1.875 366.005 2.205 ;
        RECT 365.675 0.515 366.005 0.845 ;
        RECT 365.675 -0.845 366.005 -0.515 ;
        RECT 365.68 -1.52 366 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 367.035 8.675 367.365 9.005 ;
        RECT 367.035 7.315 367.365 7.645 ;
        RECT 367.035 1.875 367.365 2.205 ;
        RECT 367.035 0.515 367.365 0.845 ;
        RECT 367.035 -0.845 367.365 -0.515 ;
        RECT 367.04 -1.52 367.36 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 368.395 8.675 368.725 9.005 ;
        RECT 368.395 7.315 368.725 7.645 ;
        RECT 368.395 1.875 368.725 2.205 ;
        RECT 368.395 0.515 368.725 0.845 ;
        RECT 368.395 -0.845 368.725 -0.515 ;
        RECT 368.4 -1.52 368.72 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 369.755 8.675 370.085 9.005 ;
        RECT 369.755 7.315 370.085 7.645 ;
        RECT 369.755 1.875 370.085 2.205 ;
        RECT 369.755 0.515 370.085 0.845 ;
        RECT 369.755 -0.845 370.085 -0.515 ;
        RECT 369.76 -1.52 370.08 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 371.115 8.675 371.445 9.005 ;
        RECT 371.115 7.315 371.445 7.645 ;
        RECT 371.115 1.875 371.445 2.205 ;
        RECT 371.115 0.515 371.445 0.845 ;
        RECT 371.115 -0.845 371.445 -0.515 ;
        RECT 371.12 -1.52 371.44 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 372.475 8.675 372.805 9.005 ;
        RECT 372.475 7.315 372.805 7.645 ;
        RECT 372.475 1.875 372.805 2.205 ;
        RECT 372.475 0.515 372.805 0.845 ;
        RECT 372.475 -0.845 372.805 -0.515 ;
        RECT 372.48 -1.52 372.8 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 373.835 8.675 374.165 9.005 ;
        RECT 373.835 7.315 374.165 7.645 ;
        RECT 373.835 1.875 374.165 2.205 ;
        RECT 373.835 0.515 374.165 0.845 ;
        RECT 373.835 -0.845 374.165 -0.515 ;
        RECT 373.84 -1.52 374.16 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 375.195 8.675 375.525 9.005 ;
        RECT 375.195 7.315 375.525 7.645 ;
        RECT 375.195 3.235 375.525 3.565 ;
        RECT 375.195 1.875 375.525 2.205 ;
        RECT 375.195 0.515 375.525 0.845 ;
        RECT 375.195 -0.845 375.525 -0.515 ;
        RECT 375.2 -1.52 375.52 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 376.555 8.675 376.885 9.005 ;
        RECT 376.555 7.315 376.885 7.645 ;
        RECT 376.555 3.235 376.885 3.565 ;
        RECT 376.555 1.875 376.885 2.205 ;
        RECT 376.555 0.515 376.885 0.845 ;
        RECT 376.555 -0.845 376.885 -0.515 ;
        RECT 376.56 -1.52 376.88 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 377.915 8.675 378.245 9.005 ;
        RECT 377.915 7.315 378.245 7.645 ;
        RECT 377.915 3.235 378.245 3.565 ;
        RECT 377.915 1.875 378.245 2.205 ;
        RECT 377.915 0.515 378.245 0.845 ;
        RECT 377.915 -0.845 378.245 -0.515 ;
        RECT 377.92 -1.52 378.24 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 379.275 8.675 379.605 9.005 ;
        RECT 379.275 7.315 379.605 7.645 ;
        RECT 379.275 1.875 379.605 2.205 ;
        RECT 379.275 0.515 379.605 0.845 ;
        RECT 379.275 -0.845 379.605 -0.515 ;
        RECT 379.28 -1.52 379.6 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 380.635 8.675 380.965 9.005 ;
        RECT 380.635 7.315 380.965 7.645 ;
        RECT 380.635 1.875 380.965 2.205 ;
        RECT 380.635 0.515 380.965 0.845 ;
        RECT 380.635 -0.845 380.965 -0.515 ;
        RECT 380.64 -1.52 380.96 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 381.995 8.675 382.325 9.005 ;
        RECT 381.995 7.315 382.325 7.645 ;
        RECT 381.995 1.875 382.325 2.205 ;
        RECT 381.995 0.515 382.325 0.845 ;
        RECT 381.995 -0.845 382.325 -0.515 ;
        RECT 382 -1.52 382.32 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 383.355 8.675 383.685 9.005 ;
        RECT 383.355 7.315 383.685 7.645 ;
        RECT 383.355 1.875 383.685 2.205 ;
        RECT 383.355 0.515 383.685 0.845 ;
        RECT 383.355 -0.845 383.685 -0.515 ;
        RECT 383.36 -1.52 383.68 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 384.715 8.675 385.045 9.005 ;
        RECT 384.715 7.315 385.045 7.645 ;
        RECT 384.715 1.875 385.045 2.205 ;
        RECT 384.715 0.515 385.045 0.845 ;
        RECT 384.715 -0.845 385.045 -0.515 ;
        RECT 384.72 -1.52 385.04 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 386.075 8.675 386.405 9.005 ;
        RECT 386.075 7.315 386.405 7.645 ;
        RECT 386.075 1.875 386.405 2.205 ;
        RECT 386.075 0.515 386.405 0.845 ;
        RECT 386.075 -0.845 386.405 -0.515 ;
        RECT 386.08 -1.52 386.4 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 387.435 8.675 387.765 9.005 ;
        RECT 387.435 7.315 387.765 7.645 ;
        RECT 387.435 3.235 387.765 3.565 ;
        RECT 387.435 1.875 387.765 2.205 ;
        RECT 387.435 0.515 387.765 0.845 ;
        RECT 387.435 -0.845 387.765 -0.515 ;
        RECT 387.44 -1.52 387.76 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 388.795 8.675 389.125 9.005 ;
        RECT 388.795 7.315 389.125 7.645 ;
        RECT 388.795 3.235 389.125 3.565 ;
        RECT 388.795 1.875 389.125 2.205 ;
        RECT 388.795 0.515 389.125 0.845 ;
        RECT 388.795 -0.845 389.125 -0.515 ;
        RECT 388.8 -1.52 389.12 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 390.155 8.675 390.485 9.005 ;
        RECT 390.155 7.315 390.485 7.645 ;
        RECT 390.155 3.235 390.485 3.565 ;
        RECT 390.155 1.875 390.485 2.205 ;
        RECT 390.155 0.515 390.485 0.845 ;
        RECT 390.155 -0.845 390.485 -0.515 ;
        RECT 390.16 -1.52 390.48 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 391.515 8.675 391.845 9.005 ;
        RECT 391.515 7.315 391.845 7.645 ;
        RECT 391.515 1.875 391.845 2.205 ;
        RECT 391.515 0.515 391.845 0.845 ;
        RECT 391.515 -0.845 391.845 -0.515 ;
        RECT 391.52 -1.52 391.84 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 392.875 8.675 393.205 9.005 ;
        RECT 392.875 7.315 393.205 7.645 ;
        RECT 392.875 1.875 393.205 2.205 ;
        RECT 392.875 0.515 393.205 0.845 ;
        RECT 392.875 -0.845 393.205 -0.515 ;
        RECT 392.88 -1.52 393.2 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 394.235 8.675 394.565 9.005 ;
        RECT 394.235 7.315 394.565 7.645 ;
        RECT 394.235 1.875 394.565 2.205 ;
        RECT 394.235 0.515 394.565 0.845 ;
        RECT 394.235 -0.845 394.565 -0.515 ;
        RECT 394.24 -1.52 394.56 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 395.595 8.675 395.925 9.005 ;
        RECT 395.595 7.315 395.925 7.645 ;
        RECT 395.595 1.875 395.925 2.205 ;
        RECT 395.595 0.515 395.925 0.845 ;
        RECT 395.595 -0.845 395.925 -0.515 ;
        RECT 395.6 -1.52 395.92 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 396.955 8.675 397.285 9.005 ;
        RECT 396.955 7.315 397.285 7.645 ;
        RECT 396.955 1.875 397.285 2.205 ;
        RECT 396.955 0.515 397.285 0.845 ;
        RECT 396.955 -0.845 397.285 -0.515 ;
        RECT 396.96 -1.52 397.28 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 398.315 8.675 398.645 9.005 ;
        RECT 398.315 7.315 398.645 7.645 ;
        RECT 398.315 1.875 398.645 2.205 ;
        RECT 398.315 0.515 398.645 0.845 ;
        RECT 398.315 -0.845 398.645 -0.515 ;
        RECT 398.32 -1.52 398.64 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 399.675 8.675 400.005 9.005 ;
        RECT 399.675 7.315 400.005 7.645 ;
        RECT 399.675 3.235 400.005 3.565 ;
        RECT 399.675 1.875 400.005 2.205 ;
        RECT 399.675 0.515 400.005 0.845 ;
        RECT 399.675 -0.845 400.005 -0.515 ;
        RECT 399.68 -1.52 400 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 401.035 8.675 401.365 9.005 ;
        RECT 401.035 7.315 401.365 7.645 ;
        RECT 401.035 3.235 401.365 3.565 ;
        RECT 401.035 1.875 401.365 2.205 ;
        RECT 401.035 0.515 401.365 0.845 ;
        RECT 401.035 -0.845 401.365 -0.515 ;
        RECT 401.04 -1.52 401.36 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 402.395 8.675 402.725 9.005 ;
        RECT 402.395 7.315 402.725 7.645 ;
        RECT 402.395 3.235 402.725 3.565 ;
        RECT 402.395 1.875 402.725 2.205 ;
        RECT 402.395 0.515 402.725 0.845 ;
        RECT 402.395 -0.845 402.725 -0.515 ;
        RECT 402.4 -1.52 402.72 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 403.755 8.675 404.085 9.005 ;
        RECT 403.755 7.315 404.085 7.645 ;
        RECT 403.755 1.875 404.085 2.205 ;
        RECT 403.755 0.515 404.085 0.845 ;
        RECT 403.755 -0.845 404.085 -0.515 ;
        RECT 403.76 -1.52 404.08 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 405.115 8.675 405.445 9.005 ;
        RECT 405.115 7.315 405.445 7.645 ;
        RECT 405.115 1.875 405.445 2.205 ;
        RECT 405.115 0.515 405.445 0.845 ;
        RECT 405.115 -0.845 405.445 -0.515 ;
        RECT 405.12 -1.52 405.44 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 406.475 8.675 406.805 9.005 ;
        RECT 406.475 7.315 406.805 7.645 ;
        RECT 406.475 1.875 406.805 2.205 ;
        RECT 406.475 0.515 406.805 0.845 ;
        RECT 406.475 -0.845 406.805 -0.515 ;
        RECT 406.48 -1.52 406.8 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 407.835 8.675 408.165 9.005 ;
        RECT 407.835 7.315 408.165 7.645 ;
        RECT 407.835 1.875 408.165 2.205 ;
        RECT 407.835 0.515 408.165 0.845 ;
        RECT 407.835 -0.845 408.165 -0.515 ;
        RECT 407.84 -1.52 408.16 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 409.195 8.675 409.525 9.005 ;
        RECT 409.195 7.315 409.525 7.645 ;
        RECT 409.195 1.875 409.525 2.205 ;
        RECT 409.195 0.515 409.525 0.845 ;
        RECT 409.195 -0.845 409.525 -0.515 ;
        RECT 409.2 -1.52 409.52 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 410.555 8.675 410.885 9.005 ;
        RECT 410.555 7.315 410.885 7.645 ;
        RECT 410.555 1.875 410.885 2.205 ;
        RECT 410.555 0.515 410.885 0.845 ;
        RECT 410.555 -0.845 410.885 -0.515 ;
        RECT 410.56 -1.52 410.88 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 411.915 8.675 412.245 9.005 ;
        RECT 411.915 7.315 412.245 7.645 ;
        RECT 411.915 3.235 412.245 3.565 ;
        RECT 411.915 1.875 412.245 2.205 ;
        RECT 411.915 0.515 412.245 0.845 ;
        RECT 411.915 -0.845 412.245 -0.515 ;
        RECT 411.92 -1.52 412.24 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 413.275 8.675 413.605 9.005 ;
        RECT 413.275 7.315 413.605 7.645 ;
        RECT 413.275 3.235 413.605 3.565 ;
        RECT 413.275 1.875 413.605 2.205 ;
        RECT 413.275 0.515 413.605 0.845 ;
        RECT 413.275 -0.845 413.605 -0.515 ;
        RECT 413.28 -1.52 413.6 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 414.635 8.675 414.965 9.005 ;
        RECT 414.635 7.315 414.965 7.645 ;
        RECT 414.635 3.235 414.965 3.565 ;
        RECT 414.635 1.875 414.965 2.205 ;
        RECT 414.635 0.515 414.965 0.845 ;
        RECT 414.635 -0.845 414.965 -0.515 ;
        RECT 414.64 -1.52 414.96 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 415.995 8.675 416.325 9.005 ;
        RECT 415.995 7.315 416.325 7.645 ;
        RECT 415.995 1.875 416.325 2.205 ;
        RECT 415.995 0.515 416.325 0.845 ;
        RECT 415.995 -0.845 416.325 -0.515 ;
        RECT 416 -1.52 416.32 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 417.355 8.675 417.685 9.005 ;
        RECT 417.355 7.315 417.685 7.645 ;
        RECT 417.355 1.875 417.685 2.205 ;
        RECT 417.355 0.515 417.685 0.845 ;
        RECT 417.355 -0.845 417.685 -0.515 ;
        RECT 417.36 -1.52 417.68 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 418.715 8.675 419.045 9.005 ;
        RECT 418.715 7.315 419.045 7.645 ;
        RECT 418.715 1.875 419.045 2.205 ;
        RECT 418.715 0.515 419.045 0.845 ;
        RECT 418.715 -0.845 419.045 -0.515 ;
        RECT 418.72 -1.52 419.04 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 420.075 8.675 420.405 9.005 ;
        RECT 420.075 7.315 420.405 7.645 ;
        RECT 420.075 1.875 420.405 2.205 ;
        RECT 420.075 0.515 420.405 0.845 ;
        RECT 420.075 -0.845 420.405 -0.515 ;
        RECT 420.08 -1.52 420.4 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 421.435 8.675 421.765 9.005 ;
        RECT 421.435 7.315 421.765 7.645 ;
        RECT 421.435 1.875 421.765 2.205 ;
        RECT 421.435 0.515 421.765 0.845 ;
        RECT 421.435 -0.845 421.765 -0.515 ;
        RECT 421.44 -1.52 421.76 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 422.795 8.675 423.125 9.005 ;
        RECT 422.795 7.315 423.125 7.645 ;
        RECT 422.795 1.875 423.125 2.205 ;
        RECT 422.795 0.515 423.125 0.845 ;
        RECT 422.795 -0.845 423.125 -0.515 ;
        RECT 422.8 -1.52 423.12 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 424.155 8.675 424.485 9.005 ;
        RECT 424.155 7.315 424.485 7.645 ;
        RECT 424.155 3.235 424.485 3.565 ;
        RECT 424.155 1.875 424.485 2.205 ;
        RECT 424.155 0.515 424.485 0.845 ;
        RECT 424.155 -0.845 424.485 -0.515 ;
        RECT 424.16 -1.52 424.48 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 425.515 8.675 425.845 9.005 ;
        RECT 425.515 7.315 425.845 7.645 ;
        RECT 425.515 3.235 425.845 3.565 ;
        RECT 425.515 1.875 425.845 2.205 ;
        RECT 425.515 0.515 425.845 0.845 ;
        RECT 425.515 -0.845 425.845 -0.515 ;
        RECT 425.52 -1.52 425.84 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 426.875 8.675 427.205 9.005 ;
        RECT 426.875 7.315 427.205 7.645 ;
        RECT 426.875 1.875 427.205 2.205 ;
        RECT 426.875 0.515 427.205 0.845 ;
        RECT 426.875 -0.845 427.205 -0.515 ;
        RECT 426.88 -1.52 427.2 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 428.235 8.675 428.565 9.005 ;
        RECT 428.235 7.315 428.565 7.645 ;
        RECT 428.235 1.875 428.565 2.205 ;
        RECT 428.235 0.515 428.565 0.845 ;
        RECT 428.235 -0.845 428.565 -0.515 ;
        RECT 428.24 -1.52 428.56 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 429.595 8.675 429.925 9.005 ;
        RECT 429.595 7.315 429.925 7.645 ;
        RECT 429.595 1.875 429.925 2.205 ;
        RECT 429.595 0.515 429.925 0.845 ;
        RECT 429.595 -0.845 429.925 -0.515 ;
        RECT 429.6 -1.52 429.92 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 430.955 8.675 431.285 9.005 ;
        RECT 430.955 7.315 431.285 7.645 ;
        RECT 430.955 1.875 431.285 2.205 ;
        RECT 430.955 0.515 431.285 0.845 ;
        RECT 430.955 -0.845 431.285 -0.515 ;
        RECT 430.96 -1.52 431.28 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 432.315 8.675 432.645 9.005 ;
        RECT 432.315 7.315 432.645 7.645 ;
        RECT 432.315 1.875 432.645 2.205 ;
        RECT 432.315 0.515 432.645 0.845 ;
        RECT 432.315 -0.845 432.645 -0.515 ;
        RECT 432.32 -1.52 432.64 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 433.675 8.675 434.005 9.005 ;
        RECT 433.675 7.315 434.005 7.645 ;
        RECT 433.675 1.875 434.005 2.205 ;
        RECT 433.675 0.515 434.005 0.845 ;
        RECT 433.675 -0.845 434.005 -0.515 ;
        RECT 433.68 -1.52 434 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 435.035 8.675 435.365 9.005 ;
        RECT 435.035 7.315 435.365 7.645 ;
        RECT 435.035 3.235 435.365 3.565 ;
        RECT 435.035 1.875 435.365 2.205 ;
        RECT 435.035 0.515 435.365 0.845 ;
        RECT 435.035 -0.845 435.365 -0.515 ;
        RECT 435.04 -1.52 435.36 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 436.395 8.675 436.725 9.005 ;
        RECT 436.395 7.315 436.725 7.645 ;
        RECT 436.395 3.235 436.725 3.565 ;
        RECT 436.395 1.875 436.725 2.205 ;
        RECT 436.395 0.515 436.725 0.845 ;
        RECT 436.395 -0.845 436.725 -0.515 ;
        RECT 436.4 -1.52 436.72 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 437.755 8.675 438.085 9.005 ;
        RECT 437.755 7.315 438.085 7.645 ;
        RECT 437.755 3.235 438.085 3.565 ;
        RECT 437.755 1.875 438.085 2.205 ;
        RECT 437.755 0.515 438.085 0.845 ;
        RECT 437.755 -0.845 438.085 -0.515 ;
        RECT 437.76 -1.52 438.08 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 439.115 8.675 439.445 9.005 ;
        RECT 439.115 7.315 439.445 7.645 ;
        RECT 439.115 1.875 439.445 2.205 ;
        RECT 439.115 0.515 439.445 0.845 ;
        RECT 439.115 -0.845 439.445 -0.515 ;
        RECT 439.12 -1.52 439.44 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 440.475 8.675 440.805 9.005 ;
        RECT 440.475 7.315 440.805 7.645 ;
        RECT 440.475 1.875 440.805 2.205 ;
        RECT 440.475 0.515 440.805 0.845 ;
        RECT 440.475 -0.845 440.805 -0.515 ;
        RECT 440.48 -1.52 440.8 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 441.835 8.675 442.165 9.005 ;
        RECT 441.835 7.315 442.165 7.645 ;
        RECT 441.835 1.875 442.165 2.205 ;
        RECT 441.835 0.515 442.165 0.845 ;
        RECT 441.835 -0.845 442.165 -0.515 ;
        RECT 441.84 -1.52 442.16 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 443.195 8.675 443.525 9.005 ;
        RECT 443.195 7.315 443.525 7.645 ;
        RECT 443.195 1.875 443.525 2.205 ;
        RECT 443.195 0.515 443.525 0.845 ;
        RECT 443.195 -0.845 443.525 -0.515 ;
        RECT 443.2 -1.52 443.52 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 444.555 8.675 444.885 9.005 ;
        RECT 444.555 7.315 444.885 7.645 ;
        RECT 444.555 1.875 444.885 2.205 ;
        RECT 444.555 0.515 444.885 0.845 ;
        RECT 444.555 -0.845 444.885 -0.515 ;
        RECT 444.56 -1.52 444.88 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 445.915 8.675 446.245 9.005 ;
        RECT 445.915 7.315 446.245 7.645 ;
        RECT 445.915 1.875 446.245 2.205 ;
        RECT 445.915 0.515 446.245 0.845 ;
        RECT 445.915 -0.845 446.245 -0.515 ;
        RECT 445.92 -1.52 446.24 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 447.275 8.675 447.605 9.005 ;
        RECT 447.275 7.315 447.605 7.645 ;
        RECT 447.275 3.235 447.605 3.565 ;
        RECT 447.275 1.875 447.605 2.205 ;
        RECT 447.275 0.515 447.605 0.845 ;
        RECT 447.275 -0.845 447.605 -0.515 ;
        RECT 447.28 -1.52 447.6 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 448.635 8.675 448.965 9.005 ;
        RECT 448.635 7.315 448.965 7.645 ;
        RECT 448.635 3.235 448.965 3.565 ;
        RECT 448.635 1.875 448.965 2.205 ;
        RECT 448.635 0.515 448.965 0.845 ;
        RECT 448.635 -0.845 448.965 -0.515 ;
        RECT 448.64 -1.52 448.96 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 449.995 8.675 450.325 9.005 ;
        RECT 449.995 7.315 450.325 7.645 ;
        RECT 449.995 3.235 450.325 3.565 ;
        RECT 449.995 1.875 450.325 2.205 ;
        RECT 449.995 0.515 450.325 0.845 ;
        RECT 449.995 -0.845 450.325 -0.515 ;
        RECT 450 -1.52 450.32 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 451.355 8.675 451.685 9.005 ;
        RECT 451.355 7.315 451.685 7.645 ;
        RECT 451.355 1.875 451.685 2.205 ;
        RECT 451.355 0.515 451.685 0.845 ;
        RECT 451.355 -0.845 451.685 -0.515 ;
        RECT 451.36 -1.52 451.68 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 452.715 8.675 453.045 9.005 ;
        RECT 452.715 7.315 453.045 7.645 ;
        RECT 452.715 1.875 453.045 2.205 ;
        RECT 452.715 0.515 453.045 0.845 ;
        RECT 452.715 -0.845 453.045 -0.515 ;
        RECT 452.72 -1.52 453.04 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 454.075 8.675 454.405 9.005 ;
        RECT 454.075 7.315 454.405 7.645 ;
        RECT 454.075 1.875 454.405 2.205 ;
        RECT 454.075 0.515 454.405 0.845 ;
        RECT 454.075 -0.845 454.405 -0.515 ;
        RECT 454.08 -1.52 454.4 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 455.435 8.675 455.765 9.005 ;
        RECT 455.435 7.315 455.765 7.645 ;
        RECT 455.435 1.875 455.765 2.205 ;
        RECT 455.435 0.515 455.765 0.845 ;
        RECT 455.435 -0.845 455.765 -0.515 ;
        RECT 455.44 -1.52 455.76 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 456.795 8.675 457.125 9.005 ;
        RECT 456.795 7.315 457.125 7.645 ;
        RECT 456.795 1.875 457.125 2.205 ;
        RECT 456.795 0.515 457.125 0.845 ;
        RECT 456.795 -0.845 457.125 -0.515 ;
        RECT 456.8 -1.52 457.12 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 458.155 8.675 458.485 9.005 ;
        RECT 458.155 7.315 458.485 7.645 ;
        RECT 458.155 1.875 458.485 2.205 ;
        RECT 458.155 0.515 458.485 0.845 ;
        RECT 458.155 -0.845 458.485 -0.515 ;
        RECT 458.16 -1.52 458.48 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 459.515 8.675 459.845 9.005 ;
        RECT 459.515 7.315 459.845 7.645 ;
        RECT 459.515 3.235 459.845 3.565 ;
        RECT 459.515 1.875 459.845 2.205 ;
        RECT 459.515 0.515 459.845 0.845 ;
        RECT 459.515 -0.845 459.845 -0.515 ;
        RECT 459.52 -1.52 459.84 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 460.875 8.675 461.205 9.005 ;
        RECT 460.875 7.315 461.205 7.645 ;
        RECT 460.875 3.235 461.205 3.565 ;
        RECT 460.875 1.875 461.205 2.205 ;
        RECT 460.875 0.515 461.205 0.845 ;
        RECT 460.875 -0.845 461.205 -0.515 ;
        RECT 460.88 -1.52 461.2 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 462.235 8.675 462.565 9.005 ;
        RECT 462.235 7.315 462.565 7.645 ;
        RECT 462.235 3.235 462.565 3.565 ;
        RECT 462.235 1.875 462.565 2.205 ;
        RECT 462.235 0.515 462.565 0.845 ;
        RECT 462.235 -0.845 462.565 -0.515 ;
        RECT 462.24 -1.52 462.56 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 463.595 8.675 463.925 9.005 ;
        RECT 463.595 7.315 463.925 7.645 ;
        RECT 463.595 1.875 463.925 2.205 ;
        RECT 463.595 0.515 463.925 0.845 ;
        RECT 463.595 -0.845 463.925 -0.515 ;
        RECT 463.6 -1.52 463.92 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 464.955 8.675 465.285 9.005 ;
        RECT 464.955 7.315 465.285 7.645 ;
        RECT 464.955 1.875 465.285 2.205 ;
        RECT 464.955 0.515 465.285 0.845 ;
        RECT 464.955 -0.845 465.285 -0.515 ;
        RECT 464.96 -1.52 465.28 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 466.315 8.675 466.645 9.005 ;
        RECT 466.315 7.315 466.645 7.645 ;
        RECT 466.315 1.875 466.645 2.205 ;
        RECT 466.315 0.515 466.645 0.845 ;
        RECT 466.315 -0.845 466.645 -0.515 ;
        RECT 466.32 -1.52 466.64 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 467.675 8.675 468.005 9.005 ;
        RECT 467.675 7.315 468.005 7.645 ;
        RECT 467.675 1.875 468.005 2.205 ;
        RECT 467.675 0.515 468.005 0.845 ;
        RECT 467.675 -0.845 468.005 -0.515 ;
        RECT 467.68 -1.52 468 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 469.035 8.675 469.365 9.005 ;
        RECT 469.035 7.315 469.365 7.645 ;
        RECT 469.035 1.875 469.365 2.205 ;
        RECT 469.035 0.515 469.365 0.845 ;
        RECT 469.035 -0.845 469.365 -0.515 ;
        RECT 469.04 -1.52 469.36 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 470.395 8.675 470.725 9.005 ;
        RECT 470.395 7.315 470.725 7.645 ;
        RECT 470.395 1.875 470.725 2.205 ;
        RECT 470.395 0.515 470.725 0.845 ;
        RECT 470.395 -0.845 470.725 -0.515 ;
        RECT 470.4 -1.52 470.72 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 471.755 8.675 472.085 9.005 ;
        RECT 471.755 7.315 472.085 7.645 ;
        RECT 471.755 3.235 472.085 3.565 ;
        RECT 471.755 1.875 472.085 2.205 ;
        RECT 471.755 0.515 472.085 0.845 ;
        RECT 471.755 -0.845 472.085 -0.515 ;
        RECT 471.76 -1.52 472.08 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 473.115 8.675 473.445 9.005 ;
        RECT 473.115 7.315 473.445 7.645 ;
        RECT 473.115 3.235 473.445 3.565 ;
        RECT 473.115 1.875 473.445 2.205 ;
        RECT 473.115 0.515 473.445 0.845 ;
        RECT 473.115 -0.845 473.445 -0.515 ;
        RECT 473.12 -1.52 473.44 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 474.475 8.675 474.805 9.005 ;
        RECT 474.475 7.315 474.805 7.645 ;
        RECT 474.475 3.235 474.805 3.565 ;
        RECT 474.475 1.875 474.805 2.205 ;
        RECT 474.475 0.515 474.805 0.845 ;
        RECT 474.475 -0.845 474.805 -0.515 ;
        RECT 474.48 -1.52 474.8 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 475.835 8.675 476.165 9.005 ;
        RECT 475.835 7.315 476.165 7.645 ;
        RECT 475.835 1.875 476.165 2.205 ;
        RECT 475.835 0.515 476.165 0.845 ;
        RECT 475.835 -0.845 476.165 -0.515 ;
        RECT 475.84 -1.52 476.16 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 477.195 8.675 477.525 9.005 ;
        RECT 477.195 7.315 477.525 7.645 ;
        RECT 477.195 1.875 477.525 2.205 ;
        RECT 477.195 0.515 477.525 0.845 ;
        RECT 477.195 -0.845 477.525 -0.515 ;
        RECT 477.2 -1.52 477.52 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 478.555 8.675 478.885 9.005 ;
        RECT 478.555 7.315 478.885 7.645 ;
        RECT 478.555 1.875 478.885 2.205 ;
        RECT 478.555 0.515 478.885 0.845 ;
        RECT 478.555 -0.845 478.885 -0.515 ;
        RECT 478.56 -1.52 478.88 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 479.915 8.675 480.245 9.005 ;
        RECT 479.915 7.315 480.245 7.645 ;
        RECT 479.915 1.875 480.245 2.205 ;
        RECT 479.915 0.515 480.245 0.845 ;
        RECT 479.915 -0.845 480.245 -0.515 ;
        RECT 479.92 -1.52 480.24 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 481.275 8.675 481.605 9.005 ;
        RECT 481.275 7.315 481.605 7.645 ;
        RECT 481.275 1.875 481.605 2.205 ;
        RECT 481.275 0.515 481.605 0.845 ;
        RECT 481.275 -0.845 481.605 -0.515 ;
        RECT 481.28 -1.52 481.6 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 482.635 8.675 482.965 9.005 ;
        RECT 482.635 7.315 482.965 7.645 ;
        RECT 482.635 1.875 482.965 2.205 ;
        RECT 482.635 0.515 482.965 0.845 ;
        RECT 482.635 -0.845 482.965 -0.515 ;
        RECT 482.64 -1.52 482.96 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 483.995 8.675 484.325 9.005 ;
        RECT 483.995 7.315 484.325 7.645 ;
        RECT 483.995 3.235 484.325 3.565 ;
        RECT 483.995 1.875 484.325 2.205 ;
        RECT 483.995 0.515 484.325 0.845 ;
        RECT 483.995 -0.845 484.325 -0.515 ;
        RECT 484 -1.52 484.32 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 485.355 8.675 485.685 9.005 ;
        RECT 485.355 7.315 485.685 7.645 ;
        RECT 485.355 3.235 485.685 3.565 ;
        RECT 485.355 1.875 485.685 2.205 ;
        RECT 485.355 0.515 485.685 0.845 ;
        RECT 485.355 -0.845 485.685 -0.515 ;
        RECT 485.36 -1.52 485.68 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 486.715 8.675 487.045 9.005 ;
        RECT 486.715 7.315 487.045 7.645 ;
        RECT 486.715 3.235 487.045 3.565 ;
        RECT 486.715 1.875 487.045 2.205 ;
        RECT 486.715 0.515 487.045 0.845 ;
        RECT 486.715 -0.845 487.045 -0.515 ;
        RECT 486.72 -1.52 487.04 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 488.075 8.675 488.405 9.005 ;
        RECT 488.075 7.315 488.405 7.645 ;
        RECT 488.075 1.875 488.405 2.205 ;
        RECT 488.075 0.515 488.405 0.845 ;
        RECT 488.075 -0.845 488.405 -0.515 ;
        RECT 488.08 -1.52 488.4 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 489.435 8.675 489.765 9.005 ;
        RECT 489.435 7.315 489.765 7.645 ;
        RECT 489.435 1.875 489.765 2.205 ;
        RECT 489.435 0.515 489.765 0.845 ;
        RECT 489.435 -0.845 489.765 -0.515 ;
        RECT 489.44 -1.52 489.76 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 490.795 8.675 491.125 9.005 ;
        RECT 490.795 7.315 491.125 7.645 ;
        RECT 490.795 1.875 491.125 2.205 ;
        RECT 490.795 0.515 491.125 0.845 ;
        RECT 490.795 -0.845 491.125 -0.515 ;
        RECT 490.8 -1.52 491.12 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 492.155 8.675 492.485 9.005 ;
        RECT 492.155 7.315 492.485 7.645 ;
        RECT 492.155 1.875 492.485 2.205 ;
        RECT 492.155 0.515 492.485 0.845 ;
        RECT 492.155 -0.845 492.485 -0.515 ;
        RECT 492.16 -1.52 492.48 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 493.515 8.675 493.845 9.005 ;
        RECT 493.515 7.315 493.845 7.645 ;
        RECT 493.515 1.875 493.845 2.205 ;
        RECT 493.515 0.515 493.845 0.845 ;
        RECT 493.515 -0.845 493.845 -0.515 ;
        RECT 493.52 -1.52 493.84 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 494.875 8.675 495.205 9.005 ;
        RECT 494.875 7.315 495.205 7.645 ;
        RECT 494.875 3.235 495.205 3.565 ;
        RECT 494.875 1.875 495.205 2.205 ;
        RECT 494.875 0.515 495.205 0.845 ;
        RECT 494.875 -0.845 495.205 -0.515 ;
        RECT 494.88 -1.52 495.2 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 496.235 8.675 496.565 9.005 ;
        RECT 496.235 7.315 496.565 7.645 ;
        RECT 496.235 3.235 496.565 3.565 ;
        RECT 496.235 1.875 496.565 2.205 ;
        RECT 496.235 0.515 496.565 0.845 ;
        RECT 496.235 -0.845 496.565 -0.515 ;
        RECT 496.24 -1.52 496.56 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 497.595 8.675 497.925 9.005 ;
        RECT 497.595 7.315 497.925 7.645 ;
        RECT 497.595 3.235 497.925 3.565 ;
        RECT 497.595 1.875 497.925 2.205 ;
        RECT 497.595 0.515 497.925 0.845 ;
        RECT 497.595 -0.845 497.925 -0.515 ;
        RECT 497.6 -1.52 497.92 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 498.955 8.675 499.285 9.005 ;
        RECT 498.955 7.315 499.285 7.645 ;
        RECT 498.955 1.875 499.285 2.205 ;
        RECT 498.955 0.515 499.285 0.845 ;
        RECT 498.955 -0.845 499.285 -0.515 ;
        RECT 498.96 -1.52 499.28 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 500.315 8.675 500.645 9.005 ;
        RECT 500.315 7.315 500.645 7.645 ;
        RECT 500.315 1.875 500.645 2.205 ;
        RECT 500.315 0.515 500.645 0.845 ;
        RECT 500.315 -0.845 500.645 -0.515 ;
        RECT 500.32 -1.52 500.64 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 501.675 8.675 502.005 9.005 ;
        RECT 501.675 7.315 502.005 7.645 ;
        RECT 501.675 1.875 502.005 2.205 ;
        RECT 501.675 0.515 502.005 0.845 ;
        RECT 501.675 -0.845 502.005 -0.515 ;
        RECT 501.68 -1.52 502 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 503.035 8.675 503.365 9.005 ;
        RECT 503.035 7.315 503.365 7.645 ;
        RECT 503.035 1.875 503.365 2.205 ;
        RECT 503.035 0.515 503.365 0.845 ;
        RECT 503.035 -0.845 503.365 -0.515 ;
        RECT 503.04 -1.52 503.36 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 504.395 8.675 504.725 9.005 ;
        RECT 504.395 7.315 504.725 7.645 ;
        RECT 504.395 1.875 504.725 2.205 ;
        RECT 504.395 0.515 504.725 0.845 ;
        RECT 504.395 -0.845 504.725 -0.515 ;
        RECT 504.4 -1.52 504.72 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 505.755 8.675 506.085 9.005 ;
        RECT 505.755 7.315 506.085 7.645 ;
        RECT 505.755 1.875 506.085 2.205 ;
        RECT 505.755 0.515 506.085 0.845 ;
        RECT 505.755 -0.845 506.085 -0.515 ;
        RECT 505.76 -1.52 506.08 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 507.115 8.675 507.445 9.005 ;
        RECT 507.115 7.315 507.445 7.645 ;
        RECT 507.115 3.235 507.445 3.565 ;
        RECT 507.115 1.875 507.445 2.205 ;
        RECT 507.115 0.515 507.445 0.845 ;
        RECT 507.115 -0.845 507.445 -0.515 ;
        RECT 507.12 -1.52 507.44 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 508.475 8.675 508.805 9.005 ;
        RECT 508.475 7.315 508.805 7.645 ;
        RECT 508.475 3.235 508.805 3.565 ;
        RECT 508.475 1.875 508.805 2.205 ;
        RECT 508.475 0.515 508.805 0.845 ;
        RECT 508.475 -0.845 508.805 -0.515 ;
        RECT 508.48 -1.52 508.8 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 509.835 8.675 510.165 9.005 ;
        RECT 509.835 7.315 510.165 7.645 ;
        RECT 509.835 3.235 510.165 3.565 ;
        RECT 509.835 1.875 510.165 2.205 ;
        RECT 509.835 0.515 510.165 0.845 ;
        RECT 509.835 -0.845 510.165 -0.515 ;
        RECT 509.84 -1.52 510.16 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 511.195 8.675 511.525 9.005 ;
        RECT 511.195 7.315 511.525 7.645 ;
        RECT 511.195 1.875 511.525 2.205 ;
        RECT 511.195 0.515 511.525 0.845 ;
        RECT 511.195 -0.845 511.525 -0.515 ;
        RECT 511.2 -1.52 511.52 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 512.555 8.675 512.885 9.005 ;
        RECT 512.555 7.315 512.885 7.645 ;
        RECT 512.555 1.875 512.885 2.205 ;
        RECT 512.555 0.515 512.885 0.845 ;
        RECT 512.555 -0.845 512.885 -0.515 ;
        RECT 512.56 -1.52 512.88 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 513.915 8.675 514.245 9.005 ;
        RECT 513.915 7.315 514.245 7.645 ;
        RECT 513.915 1.875 514.245 2.205 ;
        RECT 513.915 0.515 514.245 0.845 ;
        RECT 513.915 -0.845 514.245 -0.515 ;
        RECT 513.92 -1.52 514.24 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 515.275 8.675 515.605 9.005 ;
        RECT 515.275 7.315 515.605 7.645 ;
        RECT 515.275 1.875 515.605 2.205 ;
        RECT 515.275 0.515 515.605 0.845 ;
        RECT 515.275 -0.845 515.605 -0.515 ;
        RECT 515.28 -1.52 515.6 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 516.635 8.675 516.965 9.005 ;
        RECT 516.635 7.315 516.965 7.645 ;
        RECT 516.635 1.875 516.965 2.205 ;
        RECT 516.635 0.515 516.965 0.845 ;
        RECT 516.635 -0.845 516.965 -0.515 ;
        RECT 516.64 -1.52 516.96 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 517.995 8.675 518.325 9.005 ;
        RECT 517.995 7.315 518.325 7.645 ;
        RECT 517.995 1.875 518.325 2.205 ;
        RECT 517.995 0.515 518.325 0.845 ;
        RECT 517.995 -0.845 518.325 -0.515 ;
        RECT 518 -1.52 518.32 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 519.355 8.675 519.685 9.005 ;
        RECT 519.355 7.315 519.685 7.645 ;
        RECT 519.355 3.235 519.685 3.565 ;
        RECT 519.355 1.875 519.685 2.205 ;
        RECT 519.355 0.515 519.685 0.845 ;
        RECT 519.355 -0.845 519.685 -0.515 ;
        RECT 519.36 -1.52 519.68 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 520.715 8.675 521.045 9.005 ;
        RECT 520.715 7.315 521.045 7.645 ;
        RECT 520.715 3.235 521.045 3.565 ;
        RECT 520.715 1.875 521.045 2.205 ;
        RECT 520.715 0.515 521.045 0.845 ;
        RECT 520.715 -0.845 521.045 -0.515 ;
        RECT 520.72 -1.52 521.04 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 522.075 8.675 522.405 9.005 ;
        RECT 522.075 7.315 522.405 7.645 ;
        RECT 522.075 3.235 522.405 3.565 ;
        RECT 522.075 1.875 522.405 2.205 ;
        RECT 522.075 0.515 522.405 0.845 ;
        RECT 522.075 -0.845 522.405 -0.515 ;
        RECT 522.08 -1.52 522.4 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 523.435 8.675 523.765 9.005 ;
        RECT 523.435 7.315 523.765 7.645 ;
        RECT 523.435 1.875 523.765 2.205 ;
        RECT 523.435 0.515 523.765 0.845 ;
        RECT 523.435 -0.845 523.765 -0.515 ;
        RECT 523.44 -1.52 523.76 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 524.795 8.675 525.125 9.005 ;
        RECT 524.795 7.315 525.125 7.645 ;
        RECT 524.795 1.875 525.125 2.205 ;
        RECT 524.795 0.515 525.125 0.845 ;
        RECT 524.795 -0.845 525.125 -0.515 ;
        RECT 524.8 -1.52 525.12 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 526.155 8.675 526.485 9.005 ;
        RECT 526.155 7.315 526.485 7.645 ;
        RECT 526.155 1.875 526.485 2.205 ;
        RECT 526.155 0.515 526.485 0.845 ;
        RECT 526.155 -0.845 526.485 -0.515 ;
        RECT 526.16 -1.52 526.48 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 527.515 8.675 527.845 9.005 ;
        RECT 527.515 7.315 527.845 7.645 ;
        RECT 527.515 1.875 527.845 2.205 ;
        RECT 527.515 0.515 527.845 0.845 ;
        RECT 527.515 -0.845 527.845 -0.515 ;
        RECT 527.52 -1.52 527.84 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 528.875 8.675 529.205 9.005 ;
        RECT 528.875 7.315 529.205 7.645 ;
        RECT 528.875 1.875 529.205 2.205 ;
        RECT 528.875 0.515 529.205 0.845 ;
        RECT 528.875 -0.845 529.205 -0.515 ;
        RECT 528.88 -1.52 529.2 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 530.235 8.675 530.565 9.005 ;
        RECT 530.235 7.315 530.565 7.645 ;
        RECT 530.235 1.875 530.565 2.205 ;
        RECT 530.235 0.515 530.565 0.845 ;
        RECT 530.235 -0.845 530.565 -0.515 ;
        RECT 530.24 -1.52 530.56 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 531.595 8.675 531.925 9.005 ;
        RECT 531.595 7.315 531.925 7.645 ;
        RECT 531.595 3.235 531.925 3.565 ;
        RECT 531.595 1.875 531.925 2.205 ;
        RECT 531.595 0.515 531.925 0.845 ;
        RECT 531.595 -0.845 531.925 -0.515 ;
        RECT 531.6 -1.52 531.92 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 532.955 8.675 533.285 9.005 ;
        RECT 532.955 7.315 533.285 7.645 ;
        RECT 532.955 3.235 533.285 3.565 ;
        RECT 532.955 1.875 533.285 2.205 ;
        RECT 532.955 0.515 533.285 0.845 ;
        RECT 532.955 -0.845 533.285 -0.515 ;
        RECT 532.96 -1.52 533.28 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 534.315 8.675 534.645 9.005 ;
        RECT 534.315 7.315 534.645 7.645 ;
        RECT 534.315 3.235 534.645 3.565 ;
        RECT 534.315 1.875 534.645 2.205 ;
        RECT 534.315 0.515 534.645 0.845 ;
        RECT 534.315 -0.845 534.645 -0.515 ;
        RECT 534.32 -1.52 534.64 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 535.675 8.675 536.005 9.005 ;
        RECT 535.675 7.315 536.005 7.645 ;
        RECT 535.675 1.875 536.005 2.205 ;
        RECT 535.675 0.515 536.005 0.845 ;
        RECT 535.675 -0.845 536.005 -0.515 ;
        RECT 535.68 -1.52 536 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 537.035 8.675 537.365 9.005 ;
        RECT 537.035 7.315 537.365 7.645 ;
        RECT 537.035 1.875 537.365 2.205 ;
        RECT 537.035 0.515 537.365 0.845 ;
        RECT 537.035 -0.845 537.365 -0.515 ;
        RECT 537.04 -1.52 537.36 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 538.395 8.675 538.725 9.005 ;
        RECT 538.395 7.315 538.725 7.645 ;
        RECT 538.395 1.875 538.725 2.205 ;
        RECT 538.395 0.515 538.725 0.845 ;
        RECT 538.395 -0.845 538.725 -0.515 ;
        RECT 538.4 -1.52 538.72 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 539.755 8.675 540.085 9.005 ;
        RECT 539.755 7.315 540.085 7.645 ;
        RECT 539.755 1.875 540.085 2.205 ;
        RECT 539.755 0.515 540.085 0.845 ;
        RECT 539.755 -0.845 540.085 -0.515 ;
        RECT 539.76 -1.52 540.08 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 541.115 8.675 541.445 9.005 ;
        RECT 541.115 7.315 541.445 7.645 ;
        RECT 541.115 1.875 541.445 2.205 ;
        RECT 541.115 0.515 541.445 0.845 ;
        RECT 541.115 -0.845 541.445 -0.515 ;
        RECT 541.12 -1.52 541.44 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 542.475 8.675 542.805 9.005 ;
        RECT 542.475 7.315 542.805 7.645 ;
        RECT 542.475 1.875 542.805 2.205 ;
        RECT 542.475 0.515 542.805 0.845 ;
        RECT 542.475 -0.845 542.805 -0.515 ;
        RECT 542.48 -1.52 542.8 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 543.835 8.675 544.165 9.005 ;
        RECT 543.835 7.315 544.165 7.645 ;
        RECT 543.835 3.235 544.165 3.565 ;
        RECT 543.835 1.875 544.165 2.205 ;
        RECT 543.835 0.515 544.165 0.845 ;
        RECT 543.835 -0.845 544.165 -0.515 ;
        RECT 543.84 -1.52 544.16 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 545.195 8.675 545.525 9.005 ;
        RECT 545.195 7.315 545.525 7.645 ;
        RECT 545.195 3.235 545.525 3.565 ;
        RECT 545.195 1.875 545.525 2.205 ;
        RECT 545.195 0.515 545.525 0.845 ;
        RECT 545.195 -0.845 545.525 -0.515 ;
        RECT 545.2 -1.52 545.52 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 546.555 8.675 546.885 9.005 ;
        RECT 546.555 7.315 546.885 7.645 ;
        RECT 546.555 3.235 546.885 3.565 ;
        RECT 546.555 1.875 546.885 2.205 ;
        RECT 546.555 0.515 546.885 0.845 ;
        RECT 546.555 -0.845 546.885 -0.515 ;
        RECT 546.56 -1.52 546.88 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 547.915 8.675 548.245 9.005 ;
        RECT 547.915 7.315 548.245 7.645 ;
        RECT 547.915 1.875 548.245 2.205 ;
        RECT 547.915 0.515 548.245 0.845 ;
        RECT 547.915 -0.845 548.245 -0.515 ;
        RECT 547.92 -1.52 548.24 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 549.275 8.675 549.605 9.005 ;
        RECT 549.275 7.315 549.605 7.645 ;
        RECT 549.275 1.875 549.605 2.205 ;
        RECT 549.275 0.515 549.605 0.845 ;
        RECT 549.275 -0.845 549.605 -0.515 ;
        RECT 549.28 -1.52 549.6 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 550.635 8.675 550.965 9.005 ;
        RECT 550.635 7.315 550.965 7.645 ;
        RECT 550.635 1.875 550.965 2.205 ;
        RECT 550.635 0.515 550.965 0.845 ;
        RECT 550.635 -0.845 550.965 -0.515 ;
        RECT 550.64 -1.52 550.96 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 551.995 8.675 552.325 9.005 ;
        RECT 551.995 7.315 552.325 7.645 ;
        RECT 551.995 1.875 552.325 2.205 ;
        RECT 551.995 0.515 552.325 0.845 ;
        RECT 551.995 -0.845 552.325 -0.515 ;
        RECT 552 -1.52 552.32 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 553.355 8.675 553.685 9.005 ;
        RECT 553.355 7.315 553.685 7.645 ;
        RECT 553.355 1.875 553.685 2.205 ;
        RECT 553.355 0.515 553.685 0.845 ;
        RECT 553.355 -0.845 553.685 -0.515 ;
        RECT 553.36 -1.52 553.68 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 554.715 8.675 555.045 9.005 ;
        RECT 554.715 7.315 555.045 7.645 ;
        RECT 554.715 1.875 555.045 2.205 ;
        RECT 554.715 0.515 555.045 0.845 ;
        RECT 554.715 -0.845 555.045 -0.515 ;
        RECT 554.72 -1.52 555.04 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 556.075 0.515 556.405 0.845 ;
        RECT 556.075 -0.845 556.405 -0.515 ;
        RECT 556.08 -1.52 556.4 9.005 ;
        RECT 556.075 8.675 556.405 9.005 ;
        RECT 556.075 7.315 556.405 7.645 ;
        RECT 556.075 3.235 556.405 3.565 ;
        RECT 556.075 1.875 556.405 2.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.675 8.675 128.005 9.005 ;
        RECT 127.675 7.315 128.005 7.645 ;
        RECT 127.675 1.875 128.005 2.205 ;
        RECT 127.675 0.515 128.005 0.845 ;
        RECT 127.675 -0.845 128.005 -0.515 ;
        RECT 127.68 -1.52 128 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.035 8.675 129.365 9.005 ;
        RECT 129.035 7.315 129.365 7.645 ;
        RECT 129.035 1.875 129.365 2.205 ;
        RECT 129.035 0.515 129.365 0.845 ;
        RECT 129.035 -0.845 129.365 -0.515 ;
        RECT 129.04 -1.52 129.36 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.395 8.675 130.725 9.005 ;
        RECT 130.395 7.315 130.725 7.645 ;
        RECT 130.395 1.875 130.725 2.205 ;
        RECT 130.395 0.515 130.725 0.845 ;
        RECT 130.395 -0.845 130.725 -0.515 ;
        RECT 130.4 -1.52 130.72 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.755 8.675 132.085 9.005 ;
        RECT 131.755 7.315 132.085 7.645 ;
        RECT 131.755 1.875 132.085 2.205 ;
        RECT 131.755 0.515 132.085 0.845 ;
        RECT 131.755 -0.845 132.085 -0.515 ;
        RECT 131.76 -1.52 132.08 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.115 8.675 133.445 9.005 ;
        RECT 133.115 7.315 133.445 7.645 ;
        RECT 133.115 1.875 133.445 2.205 ;
        RECT 133.115 0.515 133.445 0.845 ;
        RECT 133.115 -0.845 133.445 -0.515 ;
        RECT 133.12 -1.52 133.44 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.475 8.675 134.805 9.005 ;
        RECT 134.475 7.315 134.805 7.645 ;
        RECT 134.475 1.875 134.805 2.205 ;
        RECT 134.475 0.515 134.805 0.845 ;
        RECT 134.475 -0.845 134.805 -0.515 ;
        RECT 134.48 -1.52 134.8 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.835 8.675 136.165 9.005 ;
        RECT 135.835 7.315 136.165 7.645 ;
        RECT 135.835 3.235 136.165 3.565 ;
        RECT 135.835 1.875 136.165 2.205 ;
        RECT 135.835 0.515 136.165 0.845 ;
        RECT 135.835 -0.845 136.165 -0.515 ;
        RECT 135.84 -1.52 136.16 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.195 8.675 137.525 9.005 ;
        RECT 137.195 7.315 137.525 7.645 ;
        RECT 137.195 3.235 137.525 3.565 ;
        RECT 137.195 1.875 137.525 2.205 ;
        RECT 137.195 0.515 137.525 0.845 ;
        RECT 137.195 -0.845 137.525 -0.515 ;
        RECT 137.2 -1.52 137.52 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 138.555 8.675 138.885 9.005 ;
        RECT 138.555 7.315 138.885 7.645 ;
        RECT 138.555 3.235 138.885 3.565 ;
        RECT 138.555 1.875 138.885 2.205 ;
        RECT 138.555 0.515 138.885 0.845 ;
        RECT 138.555 -0.845 138.885 -0.515 ;
        RECT 138.56 -1.52 138.88 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.915 8.675 140.245 9.005 ;
        RECT 139.915 7.315 140.245 7.645 ;
        RECT 139.915 1.875 140.245 2.205 ;
        RECT 139.915 0.515 140.245 0.845 ;
        RECT 139.915 -0.845 140.245 -0.515 ;
        RECT 139.92 -1.52 140.24 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.275 8.675 141.605 9.005 ;
        RECT 141.275 7.315 141.605 7.645 ;
        RECT 141.275 1.875 141.605 2.205 ;
        RECT 141.275 0.515 141.605 0.845 ;
        RECT 141.275 -0.845 141.605 -0.515 ;
        RECT 141.28 -1.52 141.6 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.635 8.675 142.965 9.005 ;
        RECT 142.635 7.315 142.965 7.645 ;
        RECT 142.635 1.875 142.965 2.205 ;
        RECT 142.635 0.515 142.965 0.845 ;
        RECT 142.635 -0.845 142.965 -0.515 ;
        RECT 142.64 -1.52 142.96 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.995 8.675 144.325 9.005 ;
        RECT 143.995 7.315 144.325 7.645 ;
        RECT 143.995 1.875 144.325 2.205 ;
        RECT 143.995 0.515 144.325 0.845 ;
        RECT 143.995 -0.845 144.325 -0.515 ;
        RECT 144 -1.52 144.32 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.355 8.675 145.685 9.005 ;
        RECT 145.355 7.315 145.685 7.645 ;
        RECT 145.355 1.875 145.685 2.205 ;
        RECT 145.355 0.515 145.685 0.845 ;
        RECT 145.355 -0.845 145.685 -0.515 ;
        RECT 145.36 -1.52 145.68 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.715 8.675 147.045 9.005 ;
        RECT 146.715 7.315 147.045 7.645 ;
        RECT 146.715 1.875 147.045 2.205 ;
        RECT 146.715 0.515 147.045 0.845 ;
        RECT 146.715 -0.845 147.045 -0.515 ;
        RECT 146.72 -1.52 147.04 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.075 8.675 148.405 9.005 ;
        RECT 148.075 7.315 148.405 7.645 ;
        RECT 148.075 3.235 148.405 3.565 ;
        RECT 148.075 1.875 148.405 2.205 ;
        RECT 148.075 0.515 148.405 0.845 ;
        RECT 148.075 -0.845 148.405 -0.515 ;
        RECT 148.08 -1.52 148.4 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.435 8.675 149.765 9.005 ;
        RECT 149.435 7.315 149.765 7.645 ;
        RECT 149.435 3.235 149.765 3.565 ;
        RECT 149.435 1.875 149.765 2.205 ;
        RECT 149.435 0.515 149.765 0.845 ;
        RECT 149.435 -0.845 149.765 -0.515 ;
        RECT 149.44 -1.52 149.76 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.795 8.675 151.125 9.005 ;
        RECT 150.795 7.315 151.125 7.645 ;
        RECT 150.795 3.235 151.125 3.565 ;
        RECT 150.795 1.875 151.125 2.205 ;
        RECT 150.795 0.515 151.125 0.845 ;
        RECT 150.795 -0.845 151.125 -0.515 ;
        RECT 150.8 -1.52 151.12 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.155 8.675 152.485 9.005 ;
        RECT 152.155 7.315 152.485 7.645 ;
        RECT 152.155 1.875 152.485 2.205 ;
        RECT 152.155 0.515 152.485 0.845 ;
        RECT 152.155 -0.845 152.485 -0.515 ;
        RECT 152.16 -1.52 152.48 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.515 8.675 153.845 9.005 ;
        RECT 153.515 7.315 153.845 7.645 ;
        RECT 153.515 1.875 153.845 2.205 ;
        RECT 153.515 0.515 153.845 0.845 ;
        RECT 153.515 -0.845 153.845 -0.515 ;
        RECT 153.52 -1.52 153.84 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.875 8.675 155.205 9.005 ;
        RECT 154.875 7.315 155.205 7.645 ;
        RECT 154.875 1.875 155.205 2.205 ;
        RECT 154.875 0.515 155.205 0.845 ;
        RECT 154.875 -0.845 155.205 -0.515 ;
        RECT 154.88 -1.52 155.2 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.235 8.675 156.565 9.005 ;
        RECT 156.235 7.315 156.565 7.645 ;
        RECT 156.235 1.875 156.565 2.205 ;
        RECT 156.235 0.515 156.565 0.845 ;
        RECT 156.235 -0.845 156.565 -0.515 ;
        RECT 156.24 -1.52 156.56 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 157.595 8.675 157.925 9.005 ;
        RECT 157.595 7.315 157.925 7.645 ;
        RECT 157.595 1.875 157.925 2.205 ;
        RECT 157.595 0.515 157.925 0.845 ;
        RECT 157.595 -0.845 157.925 -0.515 ;
        RECT 157.6 -1.52 157.92 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.955 8.675 159.285 9.005 ;
        RECT 158.955 7.315 159.285 7.645 ;
        RECT 158.955 3.235 159.285 3.565 ;
        RECT 158.955 1.875 159.285 2.205 ;
        RECT 158.955 0.515 159.285 0.845 ;
        RECT 158.955 -0.845 159.285 -0.515 ;
        RECT 158.96 -1.52 159.28 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.315 8.675 160.645 9.005 ;
        RECT 160.315 7.315 160.645 7.645 ;
        RECT 160.315 3.235 160.645 3.565 ;
        RECT 160.315 1.875 160.645 2.205 ;
        RECT 160.315 0.515 160.645 0.845 ;
        RECT 160.315 -0.845 160.645 -0.515 ;
        RECT 160.32 -1.52 160.64 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.675 8.675 162.005 9.005 ;
        RECT 161.675 7.315 162.005 7.645 ;
        RECT 161.675 3.235 162.005 3.565 ;
        RECT 161.675 1.875 162.005 2.205 ;
        RECT 161.675 0.515 162.005 0.845 ;
        RECT 161.675 -0.845 162.005 -0.515 ;
        RECT 161.68 -1.52 162 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.035 8.675 163.365 9.005 ;
        RECT 163.035 7.315 163.365 7.645 ;
        RECT 163.035 1.875 163.365 2.205 ;
        RECT 163.035 0.515 163.365 0.845 ;
        RECT 163.035 -0.845 163.365 -0.515 ;
        RECT 163.04 -1.52 163.36 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 164.395 8.675 164.725 9.005 ;
        RECT 164.395 7.315 164.725 7.645 ;
        RECT 164.395 1.875 164.725 2.205 ;
        RECT 164.395 0.515 164.725 0.845 ;
        RECT 164.395 -0.845 164.725 -0.515 ;
        RECT 164.4 -1.52 164.72 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.755 8.675 166.085 9.005 ;
        RECT 165.755 7.315 166.085 7.645 ;
        RECT 165.755 1.875 166.085 2.205 ;
        RECT 165.755 0.515 166.085 0.845 ;
        RECT 165.755 -0.845 166.085 -0.515 ;
        RECT 165.76 -1.52 166.08 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.115 8.675 167.445 9.005 ;
        RECT 167.115 7.315 167.445 7.645 ;
        RECT 167.115 1.875 167.445 2.205 ;
        RECT 167.115 0.515 167.445 0.845 ;
        RECT 167.115 -0.845 167.445 -0.515 ;
        RECT 167.12 -1.52 167.44 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 168.475 8.675 168.805 9.005 ;
        RECT 168.475 7.315 168.805 7.645 ;
        RECT 168.475 1.875 168.805 2.205 ;
        RECT 168.475 0.515 168.805 0.845 ;
        RECT 168.475 -0.845 168.805 -0.515 ;
        RECT 168.48 -1.52 168.8 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.835 8.675 170.165 9.005 ;
        RECT 169.835 7.315 170.165 7.645 ;
        RECT 169.835 1.875 170.165 2.205 ;
        RECT 169.835 0.515 170.165 0.845 ;
        RECT 169.835 -0.845 170.165 -0.515 ;
        RECT 169.84 -1.52 170.16 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.195 8.675 171.525 9.005 ;
        RECT 171.195 7.315 171.525 7.645 ;
        RECT 171.195 3.235 171.525 3.565 ;
        RECT 171.195 1.875 171.525 2.205 ;
        RECT 171.195 0.515 171.525 0.845 ;
        RECT 171.195 -0.845 171.525 -0.515 ;
        RECT 171.2 -1.52 171.52 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.555 8.675 172.885 9.005 ;
        RECT 172.555 7.315 172.885 7.645 ;
        RECT 172.555 3.235 172.885 3.565 ;
        RECT 172.555 1.875 172.885 2.205 ;
        RECT 172.555 0.515 172.885 0.845 ;
        RECT 172.555 -0.845 172.885 -0.515 ;
        RECT 172.56 -1.52 172.88 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.915 8.675 174.245 9.005 ;
        RECT 173.915 7.315 174.245 7.645 ;
        RECT 173.915 3.235 174.245 3.565 ;
        RECT 173.915 1.875 174.245 2.205 ;
        RECT 173.915 0.515 174.245 0.845 ;
        RECT 173.915 -0.845 174.245 -0.515 ;
        RECT 173.92 -1.52 174.24 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.275 8.675 175.605 9.005 ;
        RECT 175.275 7.315 175.605 7.645 ;
        RECT 175.275 1.875 175.605 2.205 ;
        RECT 175.275 0.515 175.605 0.845 ;
        RECT 175.275 -0.845 175.605 -0.515 ;
        RECT 175.28 -1.52 175.6 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 176.635 8.675 176.965 9.005 ;
        RECT 176.635 7.315 176.965 7.645 ;
        RECT 176.635 1.875 176.965 2.205 ;
        RECT 176.635 0.515 176.965 0.845 ;
        RECT 176.635 -0.845 176.965 -0.515 ;
        RECT 176.64 -1.52 176.96 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.995 8.675 178.325 9.005 ;
        RECT 177.995 7.315 178.325 7.645 ;
        RECT 177.995 1.875 178.325 2.205 ;
        RECT 177.995 0.515 178.325 0.845 ;
        RECT 177.995 -0.845 178.325 -0.515 ;
        RECT 178 -1.52 178.32 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 179.355 8.675 179.685 9.005 ;
        RECT 179.355 7.315 179.685 7.645 ;
        RECT 179.355 1.875 179.685 2.205 ;
        RECT 179.355 0.515 179.685 0.845 ;
        RECT 179.355 -0.845 179.685 -0.515 ;
        RECT 179.36 -1.52 179.68 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.715 8.675 181.045 9.005 ;
        RECT 180.715 7.315 181.045 7.645 ;
        RECT 180.715 1.875 181.045 2.205 ;
        RECT 180.715 0.515 181.045 0.845 ;
        RECT 180.715 -0.845 181.045 -0.515 ;
        RECT 180.72 -1.52 181.04 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.075 8.675 182.405 9.005 ;
        RECT 182.075 7.315 182.405 7.645 ;
        RECT 182.075 1.875 182.405 2.205 ;
        RECT 182.075 0.515 182.405 0.845 ;
        RECT 182.075 -0.845 182.405 -0.515 ;
        RECT 182.08 -1.52 182.4 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 183.435 8.675 183.765 9.005 ;
        RECT 183.435 7.315 183.765 7.645 ;
        RECT 183.435 3.235 183.765 3.565 ;
        RECT 183.435 1.875 183.765 2.205 ;
        RECT 183.435 0.515 183.765 0.845 ;
        RECT 183.435 -0.845 183.765 -0.515 ;
        RECT 183.44 -1.52 183.76 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.795 8.675 185.125 9.005 ;
        RECT 184.795 7.315 185.125 7.645 ;
        RECT 184.795 3.235 185.125 3.565 ;
        RECT 184.795 1.875 185.125 2.205 ;
        RECT 184.795 0.515 185.125 0.845 ;
        RECT 184.795 -0.845 185.125 -0.515 ;
        RECT 184.8 -1.52 185.12 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.155 8.675 186.485 9.005 ;
        RECT 186.155 7.315 186.485 7.645 ;
        RECT 186.155 3.235 186.485 3.565 ;
        RECT 186.155 1.875 186.485 2.205 ;
        RECT 186.155 0.515 186.485 0.845 ;
        RECT 186.155 -0.845 186.485 -0.515 ;
        RECT 186.16 -1.52 186.48 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 187.515 8.675 187.845 9.005 ;
        RECT 187.515 7.315 187.845 7.645 ;
        RECT 187.515 1.875 187.845 2.205 ;
        RECT 187.515 0.515 187.845 0.845 ;
        RECT 187.515 -0.845 187.845 -0.515 ;
        RECT 187.52 -1.52 187.84 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.875 8.675 189.205 9.005 ;
        RECT 188.875 7.315 189.205 7.645 ;
        RECT 188.875 1.875 189.205 2.205 ;
        RECT 188.875 0.515 189.205 0.845 ;
        RECT 188.875 -0.845 189.205 -0.515 ;
        RECT 188.88 -1.52 189.2 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.235 8.675 190.565 9.005 ;
        RECT 190.235 7.315 190.565 7.645 ;
        RECT 190.235 1.875 190.565 2.205 ;
        RECT 190.235 0.515 190.565 0.845 ;
        RECT 190.235 -0.845 190.565 -0.515 ;
        RECT 190.24 -1.52 190.56 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 191.595 8.675 191.925 9.005 ;
        RECT 191.595 7.315 191.925 7.645 ;
        RECT 191.595 1.875 191.925 2.205 ;
        RECT 191.595 0.515 191.925 0.845 ;
        RECT 191.595 -0.845 191.925 -0.515 ;
        RECT 191.6 -1.52 191.92 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.955 8.675 193.285 9.005 ;
        RECT 192.955 7.315 193.285 7.645 ;
        RECT 192.955 1.875 193.285 2.205 ;
        RECT 192.955 0.515 193.285 0.845 ;
        RECT 192.955 -0.845 193.285 -0.515 ;
        RECT 192.96 -1.52 193.28 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.315 8.675 194.645 9.005 ;
        RECT 194.315 7.315 194.645 7.645 ;
        RECT 194.315 1.875 194.645 2.205 ;
        RECT 194.315 0.515 194.645 0.845 ;
        RECT 194.315 -0.845 194.645 -0.515 ;
        RECT 194.32 -1.52 194.64 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 195.675 8.675 196.005 9.005 ;
        RECT 195.675 7.315 196.005 7.645 ;
        RECT 195.675 3.235 196.005 3.565 ;
        RECT 195.675 1.875 196.005 2.205 ;
        RECT 195.675 0.515 196.005 0.845 ;
        RECT 195.675 -0.845 196.005 -0.515 ;
        RECT 195.68 -1.52 196 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.035 8.675 197.365 9.005 ;
        RECT 197.035 7.315 197.365 7.645 ;
        RECT 197.035 3.235 197.365 3.565 ;
        RECT 197.035 1.875 197.365 2.205 ;
        RECT 197.035 0.515 197.365 0.845 ;
        RECT 197.035 -0.845 197.365 -0.515 ;
        RECT 197.04 -1.52 197.36 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.395 8.675 198.725 9.005 ;
        RECT 198.395 7.315 198.725 7.645 ;
        RECT 198.395 3.235 198.725 3.565 ;
        RECT 198.395 1.875 198.725 2.205 ;
        RECT 198.395 0.515 198.725 0.845 ;
        RECT 198.395 -0.845 198.725 -0.515 ;
        RECT 198.4 -1.52 198.72 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.755 8.675 200.085 9.005 ;
        RECT 199.755 7.315 200.085 7.645 ;
        RECT 199.755 1.875 200.085 2.205 ;
        RECT 199.755 0.515 200.085 0.845 ;
        RECT 199.755 -0.845 200.085 -0.515 ;
        RECT 199.76 -1.52 200.08 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.115 8.675 201.445 9.005 ;
        RECT 201.115 7.315 201.445 7.645 ;
        RECT 201.115 1.875 201.445 2.205 ;
        RECT 201.115 0.515 201.445 0.845 ;
        RECT 201.115 -0.845 201.445 -0.515 ;
        RECT 201.12 -1.52 201.44 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 202.475 8.675 202.805 9.005 ;
        RECT 202.475 7.315 202.805 7.645 ;
        RECT 202.475 1.875 202.805 2.205 ;
        RECT 202.475 0.515 202.805 0.845 ;
        RECT 202.475 -0.845 202.805 -0.515 ;
        RECT 202.48 -1.52 202.8 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.835 8.675 204.165 9.005 ;
        RECT 203.835 7.315 204.165 7.645 ;
        RECT 203.835 1.875 204.165 2.205 ;
        RECT 203.835 0.515 204.165 0.845 ;
        RECT 203.835 -0.845 204.165 -0.515 ;
        RECT 203.84 -1.52 204.16 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.195 8.675 205.525 9.005 ;
        RECT 205.195 7.315 205.525 7.645 ;
        RECT 205.195 1.875 205.525 2.205 ;
        RECT 205.195 0.515 205.525 0.845 ;
        RECT 205.195 -0.845 205.525 -0.515 ;
        RECT 205.2 -1.52 205.52 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 206.555 8.675 206.885 9.005 ;
        RECT 206.555 7.315 206.885 7.645 ;
        RECT 206.555 1.875 206.885 2.205 ;
        RECT 206.555 0.515 206.885 0.845 ;
        RECT 206.555 -0.845 206.885 -0.515 ;
        RECT 206.56 -1.52 206.88 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.915 8.675 208.245 9.005 ;
        RECT 207.915 7.315 208.245 7.645 ;
        RECT 207.915 3.235 208.245 3.565 ;
        RECT 207.915 1.875 208.245 2.205 ;
        RECT 207.915 0.515 208.245 0.845 ;
        RECT 207.915 -0.845 208.245 -0.515 ;
        RECT 207.92 -1.52 208.24 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.275 8.675 209.605 9.005 ;
        RECT 209.275 7.315 209.605 7.645 ;
        RECT 209.275 3.235 209.605 3.565 ;
        RECT 209.275 1.875 209.605 2.205 ;
        RECT 209.275 0.515 209.605 0.845 ;
        RECT 209.275 -0.845 209.605 -0.515 ;
        RECT 209.28 -1.52 209.6 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 210.635 8.675 210.965 9.005 ;
        RECT 210.635 7.315 210.965 7.645 ;
        RECT 210.635 3.235 210.965 3.565 ;
        RECT 210.635 1.875 210.965 2.205 ;
        RECT 210.635 0.515 210.965 0.845 ;
        RECT 210.635 -0.845 210.965 -0.515 ;
        RECT 210.64 -1.52 210.96 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 211.995 8.675 212.325 9.005 ;
        RECT 211.995 7.315 212.325 7.645 ;
        RECT 211.995 1.875 212.325 2.205 ;
        RECT 211.995 0.515 212.325 0.845 ;
        RECT 211.995 -0.845 212.325 -0.515 ;
        RECT 212 -1.52 212.32 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 213.355 8.675 213.685 9.005 ;
        RECT 213.355 7.315 213.685 7.645 ;
        RECT 213.355 1.875 213.685 2.205 ;
        RECT 213.355 0.515 213.685 0.845 ;
        RECT 213.355 -0.845 213.685 -0.515 ;
        RECT 213.36 -1.52 213.68 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.715 8.675 215.045 9.005 ;
        RECT 214.715 7.315 215.045 7.645 ;
        RECT 214.715 1.875 215.045 2.205 ;
        RECT 214.715 0.515 215.045 0.845 ;
        RECT 214.715 -0.845 215.045 -0.515 ;
        RECT 214.72 -1.52 215.04 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.075 8.675 216.405 9.005 ;
        RECT 216.075 7.315 216.405 7.645 ;
        RECT 216.075 1.875 216.405 2.205 ;
        RECT 216.075 0.515 216.405 0.845 ;
        RECT 216.075 -0.845 216.405 -0.515 ;
        RECT 216.08 -1.52 216.4 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 217.435 8.675 217.765 9.005 ;
        RECT 217.435 7.315 217.765 7.645 ;
        RECT 217.435 1.875 217.765 2.205 ;
        RECT 217.435 0.515 217.765 0.845 ;
        RECT 217.435 -0.845 217.765 -0.515 ;
        RECT 217.44 -1.52 217.76 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.795 8.675 219.125 9.005 ;
        RECT 218.795 7.315 219.125 7.645 ;
        RECT 218.795 1.875 219.125 2.205 ;
        RECT 218.795 0.515 219.125 0.845 ;
        RECT 218.795 -0.845 219.125 -0.515 ;
        RECT 218.8 -1.52 219.12 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.155 8.675 220.485 9.005 ;
        RECT 220.155 7.315 220.485 7.645 ;
        RECT 220.155 3.235 220.485 3.565 ;
        RECT 220.155 1.875 220.485 2.205 ;
        RECT 220.155 0.515 220.485 0.845 ;
        RECT 220.155 -0.845 220.485 -0.515 ;
        RECT 220.16 -1.52 220.48 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 221.515 8.675 221.845 9.005 ;
        RECT 221.515 7.315 221.845 7.645 ;
        RECT 221.515 3.235 221.845 3.565 ;
        RECT 221.515 1.875 221.845 2.205 ;
        RECT 221.515 0.515 221.845 0.845 ;
        RECT 221.515 -0.845 221.845 -0.515 ;
        RECT 221.52 -1.52 221.84 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.875 8.675 223.205 9.005 ;
        RECT 222.875 7.315 223.205 7.645 ;
        RECT 222.875 1.875 223.205 2.205 ;
        RECT 222.875 0.515 223.205 0.845 ;
        RECT 222.875 -0.845 223.205 -0.515 ;
        RECT 222.88 -1.52 223.2 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 224.235 8.675 224.565 9.005 ;
        RECT 224.235 7.315 224.565 7.645 ;
        RECT 224.235 1.875 224.565 2.205 ;
        RECT 224.235 0.515 224.565 0.845 ;
        RECT 224.235 -0.845 224.565 -0.515 ;
        RECT 224.24 -1.52 224.56 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 225.595 8.675 225.925 9.005 ;
        RECT 225.595 7.315 225.925 7.645 ;
        RECT 225.595 1.875 225.925 2.205 ;
        RECT 225.595 0.515 225.925 0.845 ;
        RECT 225.595 -0.845 225.925 -0.515 ;
        RECT 225.6 -1.52 225.92 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.955 8.675 227.285 9.005 ;
        RECT 226.955 7.315 227.285 7.645 ;
        RECT 226.955 1.875 227.285 2.205 ;
        RECT 226.955 0.515 227.285 0.845 ;
        RECT 226.955 -0.845 227.285 -0.515 ;
        RECT 226.96 -1.52 227.28 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.315 8.675 228.645 9.005 ;
        RECT 228.315 7.315 228.645 7.645 ;
        RECT 228.315 1.875 228.645 2.205 ;
        RECT 228.315 0.515 228.645 0.845 ;
        RECT 228.315 -0.845 228.645 -0.515 ;
        RECT 228.32 -1.52 228.64 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 229.675 8.675 230.005 9.005 ;
        RECT 229.675 7.315 230.005 7.645 ;
        RECT 229.675 1.875 230.005 2.205 ;
        RECT 229.675 0.515 230.005 0.845 ;
        RECT 229.675 -0.845 230.005 -0.515 ;
        RECT 229.68 -1.52 230 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 231.035 8.675 231.365 9.005 ;
        RECT 231.035 7.315 231.365 7.645 ;
        RECT 231.035 3.235 231.365 3.565 ;
        RECT 231.035 1.875 231.365 2.205 ;
        RECT 231.035 0.515 231.365 0.845 ;
        RECT 231.035 -0.845 231.365 -0.515 ;
        RECT 231.04 -1.52 231.36 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 232.395 8.675 232.725 9.005 ;
        RECT 232.395 7.315 232.725 7.645 ;
        RECT 232.395 3.235 232.725 3.565 ;
        RECT 232.395 1.875 232.725 2.205 ;
        RECT 232.395 0.515 232.725 0.845 ;
        RECT 232.395 -0.845 232.725 -0.515 ;
        RECT 232.4 -1.52 232.72 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.755 8.675 234.085 9.005 ;
        RECT 233.755 7.315 234.085 7.645 ;
        RECT 233.755 3.235 234.085 3.565 ;
        RECT 233.755 1.875 234.085 2.205 ;
        RECT 233.755 0.515 234.085 0.845 ;
        RECT 233.755 -0.845 234.085 -0.515 ;
        RECT 233.76 -1.52 234.08 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 235.115 8.675 235.445 9.005 ;
        RECT 235.115 7.315 235.445 7.645 ;
        RECT 235.115 1.875 235.445 2.205 ;
        RECT 235.115 0.515 235.445 0.845 ;
        RECT 235.115 -0.845 235.445 -0.515 ;
        RECT 235.12 -1.52 235.44 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 236.475 8.675 236.805 9.005 ;
        RECT 236.475 7.315 236.805 7.645 ;
        RECT 236.475 1.875 236.805 2.205 ;
        RECT 236.475 0.515 236.805 0.845 ;
        RECT 236.475 -0.845 236.805 -0.515 ;
        RECT 236.48 -1.52 236.8 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 237.835 8.675 238.165 9.005 ;
        RECT 237.835 7.315 238.165 7.645 ;
        RECT 237.835 1.875 238.165 2.205 ;
        RECT 237.835 0.515 238.165 0.845 ;
        RECT 237.835 -0.845 238.165 -0.515 ;
        RECT 237.84 -1.52 238.16 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.195 8.675 239.525 9.005 ;
        RECT 239.195 7.315 239.525 7.645 ;
        RECT 239.195 1.875 239.525 2.205 ;
        RECT 239.195 0.515 239.525 0.845 ;
        RECT 239.195 -0.845 239.525 -0.515 ;
        RECT 239.2 -1.52 239.52 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 240.555 8.675 240.885 9.005 ;
        RECT 240.555 7.315 240.885 7.645 ;
        RECT 240.555 1.875 240.885 2.205 ;
        RECT 240.555 0.515 240.885 0.845 ;
        RECT 240.555 -0.845 240.885 -0.515 ;
        RECT 240.56 -1.52 240.88 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 241.915 8.675 242.245 9.005 ;
        RECT 241.915 7.315 242.245 7.645 ;
        RECT 241.915 1.875 242.245 2.205 ;
        RECT 241.915 0.515 242.245 0.845 ;
        RECT 241.915 -0.845 242.245 -0.515 ;
        RECT 241.92 -1.52 242.24 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 243.275 8.675 243.605 9.005 ;
        RECT 243.275 7.315 243.605 7.645 ;
        RECT 243.275 3.235 243.605 3.565 ;
        RECT 243.275 1.875 243.605 2.205 ;
        RECT 243.275 0.515 243.605 0.845 ;
        RECT 243.275 -0.845 243.605 -0.515 ;
        RECT 243.28 -1.52 243.6 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 244.635 8.675 244.965 9.005 ;
        RECT 244.635 7.315 244.965 7.645 ;
        RECT 244.635 3.235 244.965 3.565 ;
        RECT 244.635 1.875 244.965 2.205 ;
        RECT 244.635 0.515 244.965 0.845 ;
        RECT 244.635 -0.845 244.965 -0.515 ;
        RECT 244.64 -1.52 244.96 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 245.995 8.675 246.325 9.005 ;
        RECT 245.995 7.315 246.325 7.645 ;
        RECT 245.995 3.235 246.325 3.565 ;
        RECT 245.995 1.875 246.325 2.205 ;
        RECT 245.995 0.515 246.325 0.845 ;
        RECT 245.995 -0.845 246.325 -0.515 ;
        RECT 246 -1.52 246.32 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 247.355 8.675 247.685 9.005 ;
        RECT 247.355 7.315 247.685 7.645 ;
        RECT 247.355 1.875 247.685 2.205 ;
        RECT 247.355 0.515 247.685 0.845 ;
        RECT 247.355 -0.845 247.685 -0.515 ;
        RECT 247.36 -1.52 247.68 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.715 8.675 249.045 9.005 ;
        RECT 248.715 7.315 249.045 7.645 ;
        RECT 248.715 1.875 249.045 2.205 ;
        RECT 248.715 0.515 249.045 0.845 ;
        RECT 248.715 -0.845 249.045 -0.515 ;
        RECT 248.72 -1.52 249.04 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.075 8.675 250.405 9.005 ;
        RECT 250.075 7.315 250.405 7.645 ;
        RECT 250.075 1.875 250.405 2.205 ;
        RECT 250.075 0.515 250.405 0.845 ;
        RECT 250.075 -0.845 250.405 -0.515 ;
        RECT 250.08 -1.52 250.4 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 251.435 8.675 251.765 9.005 ;
        RECT 251.435 7.315 251.765 7.645 ;
        RECT 251.435 1.875 251.765 2.205 ;
        RECT 251.435 0.515 251.765 0.845 ;
        RECT 251.435 -0.845 251.765 -0.515 ;
        RECT 251.44 -1.52 251.76 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.795 8.675 253.125 9.005 ;
        RECT 252.795 7.315 253.125 7.645 ;
        RECT 252.795 1.875 253.125 2.205 ;
        RECT 252.795 0.515 253.125 0.845 ;
        RECT 252.795 -0.845 253.125 -0.515 ;
        RECT 252.8 -1.52 253.12 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 254.155 8.675 254.485 9.005 ;
        RECT 254.155 7.315 254.485 7.645 ;
        RECT 254.155 1.875 254.485 2.205 ;
        RECT 254.155 0.515 254.485 0.845 ;
        RECT 254.155 -0.845 254.485 -0.515 ;
        RECT 254.16 -1.52 254.48 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 255.515 8.675 255.845 9.005 ;
        RECT 255.515 7.315 255.845 7.645 ;
        RECT 255.515 3.235 255.845 3.565 ;
        RECT 255.515 1.875 255.845 2.205 ;
        RECT 255.515 0.515 255.845 0.845 ;
        RECT 255.515 -0.845 255.845 -0.515 ;
        RECT 255.52 -1.52 255.84 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 256.875 8.675 257.205 9.005 ;
        RECT 256.875 7.315 257.205 7.645 ;
        RECT 256.875 3.235 257.205 3.565 ;
        RECT 256.875 1.875 257.205 2.205 ;
        RECT 256.875 0.515 257.205 0.845 ;
        RECT 256.875 -0.845 257.205 -0.515 ;
        RECT 256.88 -1.52 257.2 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.235 8.675 258.565 9.005 ;
        RECT 258.235 7.315 258.565 7.645 ;
        RECT 258.235 3.235 258.565 3.565 ;
        RECT 258.235 1.875 258.565 2.205 ;
        RECT 258.235 0.515 258.565 0.845 ;
        RECT 258.235 -0.845 258.565 -0.515 ;
        RECT 258.24 -1.52 258.56 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 259.595 8.675 259.925 9.005 ;
        RECT 259.595 7.315 259.925 7.645 ;
        RECT 259.595 1.875 259.925 2.205 ;
        RECT 259.595 0.515 259.925 0.845 ;
        RECT 259.595 -0.845 259.925 -0.515 ;
        RECT 259.6 -1.52 259.92 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.955 8.675 261.285 9.005 ;
        RECT 260.955 7.315 261.285 7.645 ;
        RECT 260.955 1.875 261.285 2.205 ;
        RECT 260.955 0.515 261.285 0.845 ;
        RECT 260.955 -0.845 261.285 -0.515 ;
        RECT 260.96 -1.52 261.28 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.315 8.675 262.645 9.005 ;
        RECT 262.315 7.315 262.645 7.645 ;
        RECT 262.315 1.875 262.645 2.205 ;
        RECT 262.315 0.515 262.645 0.845 ;
        RECT 262.315 -0.845 262.645 -0.515 ;
        RECT 262.32 -1.52 262.64 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 263.675 8.675 264.005 9.005 ;
        RECT 263.675 7.315 264.005 7.645 ;
        RECT 263.675 1.875 264.005 2.205 ;
        RECT 263.675 0.515 264.005 0.845 ;
        RECT 263.675 -0.845 264.005 -0.515 ;
        RECT 263.68 -1.52 264 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 265.035 8.675 265.365 9.005 ;
        RECT 265.035 7.315 265.365 7.645 ;
        RECT 265.035 1.875 265.365 2.205 ;
        RECT 265.035 0.515 265.365 0.845 ;
        RECT 265.035 -0.845 265.365 -0.515 ;
        RECT 265.04 -1.52 265.36 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 266.395 8.675 266.725 9.005 ;
        RECT 266.395 7.315 266.725 7.645 ;
        RECT 266.395 1.875 266.725 2.205 ;
        RECT 266.395 0.515 266.725 0.845 ;
        RECT 266.395 -0.845 266.725 -0.515 ;
        RECT 266.4 -1.52 266.72 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 267.755 8.675 268.085 9.005 ;
        RECT 267.755 7.315 268.085 7.645 ;
        RECT 267.755 3.235 268.085 3.565 ;
        RECT 267.755 1.875 268.085 2.205 ;
        RECT 267.755 0.515 268.085 0.845 ;
        RECT 267.755 -0.845 268.085 -0.515 ;
        RECT 267.76 -1.52 268.08 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.115 8.675 269.445 9.005 ;
        RECT 269.115 7.315 269.445 7.645 ;
        RECT 269.115 3.235 269.445 3.565 ;
        RECT 269.115 1.875 269.445 2.205 ;
        RECT 269.115 0.515 269.445 0.845 ;
        RECT 269.115 -0.845 269.445 -0.515 ;
        RECT 269.12 -1.52 269.44 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 270.475 8.675 270.805 9.005 ;
        RECT 270.475 7.315 270.805 7.645 ;
        RECT 270.475 3.235 270.805 3.565 ;
        RECT 270.475 1.875 270.805 2.205 ;
        RECT 270.475 0.515 270.805 0.845 ;
        RECT 270.475 -0.845 270.805 -0.515 ;
        RECT 270.48 -1.52 270.8 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.835 8.675 272.165 9.005 ;
        RECT 271.835 7.315 272.165 7.645 ;
        RECT 271.835 1.875 272.165 2.205 ;
        RECT 271.835 0.515 272.165 0.845 ;
        RECT 271.835 -0.845 272.165 -0.515 ;
        RECT 271.84 -1.52 272.16 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.195 8.675 273.525 9.005 ;
        RECT 273.195 7.315 273.525 7.645 ;
        RECT 273.195 1.875 273.525 2.205 ;
        RECT 273.195 0.515 273.525 0.845 ;
        RECT 273.195 -0.845 273.525 -0.515 ;
        RECT 273.2 -1.52 273.52 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 274.555 8.675 274.885 9.005 ;
        RECT 274.555 7.315 274.885 7.645 ;
        RECT 274.555 1.875 274.885 2.205 ;
        RECT 274.555 0.515 274.885 0.845 ;
        RECT 274.555 -0.845 274.885 -0.515 ;
        RECT 274.56 -1.52 274.88 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.915 8.675 276.245 9.005 ;
        RECT 275.915 7.315 276.245 7.645 ;
        RECT 275.915 1.875 276.245 2.205 ;
        RECT 275.915 0.515 276.245 0.845 ;
        RECT 275.915 -0.845 276.245 -0.515 ;
        RECT 275.92 -1.52 276.24 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 277.275 8.675 277.605 9.005 ;
        RECT 277.275 7.315 277.605 7.645 ;
        RECT 277.275 1.875 277.605 2.205 ;
        RECT 277.275 0.515 277.605 0.845 ;
        RECT 277.275 -0.845 277.605 -0.515 ;
        RECT 277.28 -1.52 277.6 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 278.635 8.675 278.965 9.005 ;
        RECT 278.635 7.315 278.965 7.645 ;
        RECT 278.635 1.875 278.965 2.205 ;
        RECT 278.635 0.515 278.965 0.845 ;
        RECT 278.635 -0.845 278.965 -0.515 ;
        RECT 278.64 -1.52 278.96 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.995 8.675 280.325 9.005 ;
        RECT 279.995 7.315 280.325 7.645 ;
        RECT 279.995 3.235 280.325 3.565 ;
        RECT 279.995 1.875 280.325 2.205 ;
        RECT 279.995 0.515 280.325 0.845 ;
        RECT 279.995 -0.845 280.325 -0.515 ;
        RECT 280 -1.52 280.32 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 281.355 8.675 281.685 9.005 ;
        RECT 281.355 7.315 281.685 7.645 ;
        RECT 281.355 3.235 281.685 3.565 ;
        RECT 281.355 1.875 281.685 2.205 ;
        RECT 281.355 0.515 281.685 0.845 ;
        RECT 281.355 -0.845 281.685 -0.515 ;
        RECT 281.36 -1.52 281.68 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.715 8.675 283.045 9.005 ;
        RECT 282.715 7.315 283.045 7.645 ;
        RECT 282.715 3.235 283.045 3.565 ;
        RECT 282.715 1.875 283.045 2.205 ;
        RECT 282.715 0.515 283.045 0.845 ;
        RECT 282.715 -0.845 283.045 -0.515 ;
        RECT 282.72 -1.52 283.04 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 284.075 8.675 284.405 9.005 ;
        RECT 284.075 7.315 284.405 7.645 ;
        RECT 284.075 1.875 284.405 2.205 ;
        RECT 284.075 0.515 284.405 0.845 ;
        RECT 284.075 -0.845 284.405 -0.515 ;
        RECT 284.08 -1.52 284.4 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 285.435 8.675 285.765 9.005 ;
        RECT 285.435 7.315 285.765 7.645 ;
        RECT 285.435 1.875 285.765 2.205 ;
        RECT 285.435 0.515 285.765 0.845 ;
        RECT 285.435 -0.845 285.765 -0.515 ;
        RECT 285.44 -1.52 285.76 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.795 8.675 287.125 9.005 ;
        RECT 286.795 7.315 287.125 7.645 ;
        RECT 286.795 1.875 287.125 2.205 ;
        RECT 286.795 0.515 287.125 0.845 ;
        RECT 286.795 -0.845 287.125 -0.515 ;
        RECT 286.8 -1.52 287.12 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.155 8.675 288.485 9.005 ;
        RECT 288.155 7.315 288.485 7.645 ;
        RECT 288.155 1.875 288.485 2.205 ;
        RECT 288.155 0.515 288.485 0.845 ;
        RECT 288.155 -0.845 288.485 -0.515 ;
        RECT 288.16 -1.52 288.48 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 289.515 8.675 289.845 9.005 ;
        RECT 289.515 7.315 289.845 7.645 ;
        RECT 289.515 1.875 289.845 2.205 ;
        RECT 289.515 0.515 289.845 0.845 ;
        RECT 289.515 -0.845 289.845 -0.515 ;
        RECT 289.52 -1.52 289.84 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.875 8.675 291.205 9.005 ;
        RECT 290.875 7.315 291.205 7.645 ;
        RECT 290.875 3.235 291.205 3.565 ;
        RECT 290.875 1.875 291.205 2.205 ;
        RECT 290.875 0.515 291.205 0.845 ;
        RECT 290.875 -0.845 291.205 -0.515 ;
        RECT 290.88 -1.52 291.2 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.235 8.675 292.565 9.005 ;
        RECT 292.235 7.315 292.565 7.645 ;
        RECT 292.235 3.235 292.565 3.565 ;
        RECT 292.235 1.875 292.565 2.205 ;
        RECT 292.235 0.515 292.565 0.845 ;
        RECT 292.235 -0.845 292.565 -0.515 ;
        RECT 292.24 -1.52 292.56 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 293.595 8.675 293.925 9.005 ;
        RECT 293.595 7.315 293.925 7.645 ;
        RECT 293.595 3.235 293.925 3.565 ;
        RECT 293.595 1.875 293.925 2.205 ;
        RECT 293.595 0.515 293.925 0.845 ;
        RECT 293.595 -0.845 293.925 -0.515 ;
        RECT 293.6 -1.52 293.92 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.955 8.675 295.285 9.005 ;
        RECT 294.955 7.315 295.285 7.645 ;
        RECT 294.955 1.875 295.285 2.205 ;
        RECT 294.955 0.515 295.285 0.845 ;
        RECT 294.955 -0.845 295.285 -0.515 ;
        RECT 294.96 -1.52 295.28 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 296.315 8.675 296.645 9.005 ;
        RECT 296.315 7.315 296.645 7.645 ;
        RECT 296.315 1.875 296.645 2.205 ;
        RECT 296.315 0.515 296.645 0.845 ;
        RECT 296.315 -0.845 296.645 -0.515 ;
        RECT 296.32 -1.52 296.64 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 297.675 8.675 298.005 9.005 ;
        RECT 297.675 7.315 298.005 7.645 ;
        RECT 297.675 1.875 298.005 2.205 ;
        RECT 297.675 0.515 298.005 0.845 ;
        RECT 297.675 -0.845 298.005 -0.515 ;
        RECT 297.68 -1.52 298 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 299.035 8.675 299.365 9.005 ;
        RECT 299.035 7.315 299.365 7.645 ;
        RECT 299.035 1.875 299.365 2.205 ;
        RECT 299.035 0.515 299.365 0.845 ;
        RECT 299.035 -0.845 299.365 -0.515 ;
        RECT 299.04 -1.52 299.36 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 300.395 8.675 300.725 9.005 ;
        RECT 300.395 7.315 300.725 7.645 ;
        RECT 300.395 1.875 300.725 2.205 ;
        RECT 300.395 0.515 300.725 0.845 ;
        RECT 300.395 -0.845 300.725 -0.515 ;
        RECT 300.4 -1.52 300.72 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.755 8.675 302.085 9.005 ;
        RECT 301.755 7.315 302.085 7.645 ;
        RECT 301.755 1.875 302.085 2.205 ;
        RECT 301.755 0.515 302.085 0.845 ;
        RECT 301.755 -0.845 302.085 -0.515 ;
        RECT 301.76 -1.52 302.08 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.115 8.675 303.445 9.005 ;
        RECT 303.115 7.315 303.445 7.645 ;
        RECT 303.115 3.235 303.445 3.565 ;
        RECT 303.115 1.875 303.445 2.205 ;
        RECT 303.115 0.515 303.445 0.845 ;
        RECT 303.115 -0.845 303.445 -0.515 ;
        RECT 303.12 -1.52 303.44 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 304.475 8.675 304.805 9.005 ;
        RECT 304.475 7.315 304.805 7.645 ;
        RECT 304.475 3.235 304.805 3.565 ;
        RECT 304.475 1.875 304.805 2.205 ;
        RECT 304.475 0.515 304.805 0.845 ;
        RECT 304.475 -0.845 304.805 -0.515 ;
        RECT 304.48 -1.52 304.8 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.835 8.675 306.165 9.005 ;
        RECT 305.835 7.315 306.165 7.645 ;
        RECT 305.835 3.235 306.165 3.565 ;
        RECT 305.835 1.875 306.165 2.205 ;
        RECT 305.835 0.515 306.165 0.845 ;
        RECT 305.835 -0.845 306.165 -0.515 ;
        RECT 305.84 -1.52 306.16 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.195 8.675 307.525 9.005 ;
        RECT 307.195 7.315 307.525 7.645 ;
        RECT 307.195 1.875 307.525 2.205 ;
        RECT 307.195 0.515 307.525 0.845 ;
        RECT 307.195 -0.845 307.525 -0.515 ;
        RECT 307.2 -1.52 307.52 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 308.555 8.675 308.885 9.005 ;
        RECT 308.555 7.315 308.885 7.645 ;
        RECT 308.555 1.875 308.885 2.205 ;
        RECT 308.555 0.515 308.885 0.845 ;
        RECT 308.555 -0.845 308.885 -0.515 ;
        RECT 308.56 -1.52 308.88 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.915 8.675 310.245 9.005 ;
        RECT 309.915 7.315 310.245 7.645 ;
        RECT 309.915 1.875 310.245 2.205 ;
        RECT 309.915 0.515 310.245 0.845 ;
        RECT 309.915 -0.845 310.245 -0.515 ;
        RECT 309.92 -1.52 310.24 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 311.275 8.675 311.605 9.005 ;
        RECT 311.275 7.315 311.605 7.645 ;
        RECT 311.275 1.875 311.605 2.205 ;
        RECT 311.275 0.515 311.605 0.845 ;
        RECT 311.275 -0.845 311.605 -0.515 ;
        RECT 311.28 -1.52 311.6 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 312.635 8.675 312.965 9.005 ;
        RECT 312.635 7.315 312.965 7.645 ;
        RECT 312.635 1.875 312.965 2.205 ;
        RECT 312.635 0.515 312.965 0.845 ;
        RECT 312.635 -0.845 312.965 -0.515 ;
        RECT 312.64 -1.52 312.96 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.995 8.675 314.325 9.005 ;
        RECT 313.995 7.315 314.325 7.645 ;
        RECT 313.995 1.875 314.325 2.205 ;
        RECT 313.995 0.515 314.325 0.845 ;
        RECT 313.995 -0.845 314.325 -0.515 ;
        RECT 314 -1.52 314.32 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 315.355 8.675 315.685 9.005 ;
        RECT 315.355 7.315 315.685 7.645 ;
        RECT 315.355 3.235 315.685 3.565 ;
        RECT 315.355 1.875 315.685 2.205 ;
        RECT 315.355 0.515 315.685 0.845 ;
        RECT 315.355 -0.845 315.685 -0.515 ;
        RECT 315.36 -1.52 315.68 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 316.715 8.675 317.045 9.005 ;
        RECT 316.715 7.315 317.045 7.645 ;
        RECT 316.715 3.235 317.045 3.565 ;
        RECT 316.715 1.875 317.045 2.205 ;
        RECT 316.715 0.515 317.045 0.845 ;
        RECT 316.715 -0.845 317.045 -0.515 ;
        RECT 316.72 -1.52 317.04 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.075 8.675 318.405 9.005 ;
        RECT 318.075 7.315 318.405 7.645 ;
        RECT 318.075 3.235 318.405 3.565 ;
        RECT 318.075 1.875 318.405 2.205 ;
        RECT 318.075 0.515 318.405 0.845 ;
        RECT 318.075 -0.845 318.405 -0.515 ;
        RECT 318.08 -1.52 318.4 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 319.435 8.675 319.765 9.005 ;
        RECT 319.435 7.315 319.765 7.645 ;
        RECT 319.435 1.875 319.765 2.205 ;
        RECT 319.435 0.515 319.765 0.845 ;
        RECT 319.435 -0.845 319.765 -0.515 ;
        RECT 319.44 -1.52 319.76 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 320.795 8.675 321.125 9.005 ;
        RECT 320.795 7.315 321.125 7.645 ;
        RECT 320.795 1.875 321.125 2.205 ;
        RECT 320.795 0.515 321.125 0.845 ;
        RECT 320.795 -0.845 321.125 -0.515 ;
        RECT 320.8 -1.52 321.12 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 322.155 8.675 322.485 9.005 ;
        RECT 322.155 7.315 322.485 7.645 ;
        RECT 322.155 1.875 322.485 2.205 ;
        RECT 322.155 0.515 322.485 0.845 ;
        RECT 322.155 -0.845 322.485 -0.515 ;
        RECT 322.16 -1.52 322.48 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 323.515 8.675 323.845 9.005 ;
        RECT 323.515 7.315 323.845 7.645 ;
        RECT 323.515 1.875 323.845 2.205 ;
        RECT 323.515 0.515 323.845 0.845 ;
        RECT 323.515 -0.845 323.845 -0.515 ;
        RECT 323.52 -1.52 323.84 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.875 8.675 325.205 9.005 ;
        RECT 324.875 7.315 325.205 7.645 ;
        RECT 324.875 1.875 325.205 2.205 ;
        RECT 324.875 0.515 325.205 0.845 ;
        RECT 324.875 -0.845 325.205 -0.515 ;
        RECT 324.88 -1.52 325.2 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 326.235 8.675 326.565 9.005 ;
        RECT 326.235 7.315 326.565 7.645 ;
        RECT 326.235 1.875 326.565 2.205 ;
        RECT 326.235 0.515 326.565 0.845 ;
        RECT 326.235 -0.845 326.565 -0.515 ;
        RECT 326.24 -1.52 326.56 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 327.595 8.675 327.925 9.005 ;
        RECT 327.595 7.315 327.925 7.645 ;
        RECT 327.595 3.235 327.925 3.565 ;
        RECT 327.595 1.875 327.925 2.205 ;
        RECT 327.595 0.515 327.925 0.845 ;
        RECT 327.595 -0.845 327.925 -0.515 ;
        RECT 327.6 -1.52 327.92 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 328.955 8.675 329.285 9.005 ;
        RECT 328.955 7.315 329.285 7.645 ;
        RECT 328.955 3.235 329.285 3.565 ;
        RECT 328.955 1.875 329.285 2.205 ;
        RECT 328.955 0.515 329.285 0.845 ;
        RECT 328.955 -0.845 329.285 -0.515 ;
        RECT 328.96 -1.52 329.28 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.315 8.675 330.645 9.005 ;
        RECT 330.315 7.315 330.645 7.645 ;
        RECT 330.315 3.235 330.645 3.565 ;
        RECT 330.315 1.875 330.645 2.205 ;
        RECT 330.315 0.515 330.645 0.845 ;
        RECT 330.315 -0.845 330.645 -0.515 ;
        RECT 330.32 -1.52 330.64 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 331.675 8.675 332.005 9.005 ;
        RECT 331.675 7.315 332.005 7.645 ;
        RECT 331.675 1.875 332.005 2.205 ;
        RECT 331.675 0.515 332.005 0.845 ;
        RECT 331.675 -0.845 332.005 -0.515 ;
        RECT 331.68 -1.52 332 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 333.035 8.675 333.365 9.005 ;
        RECT 333.035 7.315 333.365 7.645 ;
        RECT 333.035 1.875 333.365 2.205 ;
        RECT 333.035 0.515 333.365 0.845 ;
        RECT 333.035 -0.845 333.365 -0.515 ;
        RECT 333.04 -1.52 333.36 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 334.395 8.675 334.725 9.005 ;
        RECT 334.395 7.315 334.725 7.645 ;
        RECT 334.395 1.875 334.725 2.205 ;
        RECT 334.395 0.515 334.725 0.845 ;
        RECT 334.395 -0.845 334.725 -0.515 ;
        RECT 334.4 -1.52 334.72 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.755 8.675 336.085 9.005 ;
        RECT 335.755 7.315 336.085 7.645 ;
        RECT 335.755 1.875 336.085 2.205 ;
        RECT 335.755 0.515 336.085 0.845 ;
        RECT 335.755 -0.845 336.085 -0.515 ;
        RECT 335.76 -1.52 336.08 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 337.115 8.675 337.445 9.005 ;
        RECT 337.115 7.315 337.445 7.645 ;
        RECT 337.115 1.875 337.445 2.205 ;
        RECT 337.115 0.515 337.445 0.845 ;
        RECT 337.115 -0.845 337.445 -0.515 ;
        RECT 337.12 -1.52 337.44 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 338.475 8.675 338.805 9.005 ;
        RECT 338.475 7.315 338.805 7.645 ;
        RECT 338.475 1.875 338.805 2.205 ;
        RECT 338.475 0.515 338.805 0.845 ;
        RECT 338.475 -0.845 338.805 -0.515 ;
        RECT 338.48 -1.52 338.8 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 339.835 8.675 340.165 9.005 ;
        RECT 339.835 7.315 340.165 7.645 ;
        RECT 339.835 3.235 340.165 3.565 ;
        RECT 339.835 1.875 340.165 2.205 ;
        RECT 339.835 0.515 340.165 0.845 ;
        RECT 339.835 -0.845 340.165 -0.515 ;
        RECT 339.84 -1.52 340.16 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 341.195 0.515 341.525 0.845 ;
        RECT 341.195 -0.845 341.525 -0.515 ;
        RECT 341.2 -1.52 341.52 9.005 ;
        RECT 341.195 8.675 341.525 9.005 ;
        RECT 341.195 7.315 341.525 7.645 ;
        RECT 341.195 3.235 341.525 3.565 ;
        RECT 341.195 1.875 341.525 2.205 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.525 8.675 -1.195 9.005 ;
        RECT -1.525 7.315 -1.195 7.645 ;
        RECT -1.525 5.955 -1.195 6.285 ;
        RECT -1.525 4.595 -1.195 4.925 ;
        RECT -1.525 3.235 -1.195 3.565 ;
        RECT -1.525 1.875 -1.195 2.205 ;
        RECT -1.525 0.515 -1.195 0.845 ;
        RECT -1.525 -0.845 -1.195 -0.515 ;
        RECT -1.52 -1.52 -1.2 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.165 8.675 0.165 9.005 ;
        RECT -0.165 7.315 0.165 7.645 ;
        RECT -0.165 4.595 0.165 4.925 ;
        RECT -0.165 3.235 0.165 3.565 ;
        RECT -0.165 1.875 0.165 2.205 ;
        RECT -0.165 0.515 0.165 0.845 ;
        RECT -0.165 -0.845 0.165 -0.515 ;
        RECT -0.16 -1.52 0.16 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.195 8.675 1.525 9.005 ;
        RECT 1.195 7.315 1.525 7.645 ;
        RECT 1.195 3.235 1.525 3.565 ;
        RECT 1.195 1.875 1.525 2.205 ;
        RECT 1.195 0.515 1.525 0.845 ;
        RECT 1.195 -0.845 1.525 -0.515 ;
        RECT 1.2 -1.52 1.52 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 8.675 2.885 9.005 ;
        RECT 2.555 7.315 2.885 7.645 ;
        RECT 2.555 3.235 2.885 3.565 ;
        RECT 2.555 1.875 2.885 2.205 ;
        RECT 2.555 0.515 2.885 0.845 ;
        RECT 2.555 -0.845 2.885 -0.515 ;
        RECT 2.56 -1.52 2.88 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.915 8.675 4.245 9.005 ;
        RECT 3.915 7.315 4.245 7.645 ;
        RECT 3.915 3.235 4.245 3.565 ;
        RECT 3.915 1.875 4.245 2.205 ;
        RECT 3.915 0.515 4.245 0.845 ;
        RECT 3.915 -0.845 4.245 -0.515 ;
        RECT 3.92 -1.52 4.24 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.275 8.675 5.605 9.005 ;
        RECT 5.275 7.315 5.605 7.645 ;
        RECT 5.275 3.235 5.605 3.565 ;
        RECT 5.275 1.875 5.605 2.205 ;
        RECT 5.275 0.515 5.605 0.845 ;
        RECT 5.275 -0.845 5.605 -0.515 ;
        RECT 5.28 -1.52 5.6 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 8.675 6.965 9.005 ;
        RECT 6.635 7.315 6.965 7.645 ;
        RECT 6.635 3.235 6.965 3.565 ;
        RECT 6.635 1.875 6.965 2.205 ;
        RECT 6.635 0.515 6.965 0.845 ;
        RECT 6.635 -0.845 6.965 -0.515 ;
        RECT 6.64 -1.52 6.96 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.995 8.675 8.325 9.005 ;
        RECT 7.995 7.315 8.325 7.645 ;
        RECT 7.995 1.875 8.325 2.205 ;
        RECT 7.995 0.515 8.325 0.845 ;
        RECT 7.995 -0.845 8.325 -0.515 ;
        RECT 8 -1.52 8.32 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 8.675 9.685 9.005 ;
        RECT 9.355 7.315 9.685 7.645 ;
        RECT 9.355 1.875 9.685 2.205 ;
        RECT 9.355 0.515 9.685 0.845 ;
        RECT 9.355 -0.845 9.685 -0.515 ;
        RECT 9.36 -1.52 9.68 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.715 8.675 11.045 9.005 ;
        RECT 10.715 7.315 11.045 7.645 ;
        RECT 10.715 1.875 11.045 2.205 ;
        RECT 10.715 0.515 11.045 0.845 ;
        RECT 10.715 -0.845 11.045 -0.515 ;
        RECT 10.72 -1.52 11.04 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.075 8.675 12.405 9.005 ;
        RECT 12.075 7.315 12.405 7.645 ;
        RECT 12.075 1.875 12.405 2.205 ;
        RECT 12.075 0.515 12.405 0.845 ;
        RECT 12.075 -0.845 12.405 -0.515 ;
        RECT 12.08 -1.52 12.4 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.435 8.675 13.765 9.005 ;
        RECT 13.435 7.315 13.765 7.645 ;
        RECT 13.435 1.875 13.765 2.205 ;
        RECT 13.435 0.515 13.765 0.845 ;
        RECT 13.435 -0.845 13.765 -0.515 ;
        RECT 13.44 -1.52 13.76 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.795 8.675 15.125 9.005 ;
        RECT 14.795 7.315 15.125 7.645 ;
        RECT 14.795 1.875 15.125 2.205 ;
        RECT 14.795 0.515 15.125 0.845 ;
        RECT 14.795 -0.845 15.125 -0.515 ;
        RECT 14.8 -1.52 15.12 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.155 8.675 16.485 9.005 ;
        RECT 16.155 7.315 16.485 7.645 ;
        RECT 16.155 3.235 16.485 3.565 ;
        RECT 16.155 1.875 16.485 2.205 ;
        RECT 16.155 0.515 16.485 0.845 ;
        RECT 16.155 -0.845 16.485 -0.515 ;
        RECT 16.16 -1.52 16.48 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.515 8.675 17.845 9.005 ;
        RECT 17.515 7.315 17.845 7.645 ;
        RECT 17.515 3.235 17.845 3.565 ;
        RECT 17.515 1.875 17.845 2.205 ;
        RECT 17.515 0.515 17.845 0.845 ;
        RECT 17.515 -0.845 17.845 -0.515 ;
        RECT 17.52 -1.52 17.84 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.875 8.675 19.205 9.005 ;
        RECT 18.875 7.315 19.205 7.645 ;
        RECT 18.875 1.875 19.205 2.205 ;
        RECT 18.875 0.515 19.205 0.845 ;
        RECT 18.875 -0.845 19.205 -0.515 ;
        RECT 18.88 -1.52 19.2 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.235 8.675 20.565 9.005 ;
        RECT 20.235 7.315 20.565 7.645 ;
        RECT 20.235 1.875 20.565 2.205 ;
        RECT 20.235 0.515 20.565 0.845 ;
        RECT 20.235 -0.845 20.565 -0.515 ;
        RECT 20.24 -1.52 20.56 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.595 8.675 21.925 9.005 ;
        RECT 21.595 7.315 21.925 7.645 ;
        RECT 21.595 1.875 21.925 2.205 ;
        RECT 21.595 0.515 21.925 0.845 ;
        RECT 21.595 -0.845 21.925 -0.515 ;
        RECT 21.6 -1.52 21.92 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.955 8.675 23.285 9.005 ;
        RECT 22.955 7.315 23.285 7.645 ;
        RECT 22.955 1.875 23.285 2.205 ;
        RECT 22.955 0.515 23.285 0.845 ;
        RECT 22.955 -0.845 23.285 -0.515 ;
        RECT 22.96 -1.52 23.28 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.315 8.675 24.645 9.005 ;
        RECT 24.315 7.315 24.645 7.645 ;
        RECT 24.315 1.875 24.645 2.205 ;
        RECT 24.315 0.515 24.645 0.845 ;
        RECT 24.315 -0.845 24.645 -0.515 ;
        RECT 24.32 -1.52 24.64 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.675 8.675 26.005 9.005 ;
        RECT 25.675 7.315 26.005 7.645 ;
        RECT 25.675 1.875 26.005 2.205 ;
        RECT 25.675 0.515 26.005 0.845 ;
        RECT 25.675 -0.845 26.005 -0.515 ;
        RECT 25.68 -1.52 26 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.035 8.675 27.365 9.005 ;
        RECT 27.035 7.315 27.365 7.645 ;
        RECT 27.035 3.235 27.365 3.565 ;
        RECT 27.035 1.875 27.365 2.205 ;
        RECT 27.035 0.515 27.365 0.845 ;
        RECT 27.035 -0.845 27.365 -0.515 ;
        RECT 27.04 -1.52 27.36 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.395 8.675 28.725 9.005 ;
        RECT 28.395 7.315 28.725 7.645 ;
        RECT 28.395 3.235 28.725 3.565 ;
        RECT 28.395 1.875 28.725 2.205 ;
        RECT 28.395 0.515 28.725 0.845 ;
        RECT 28.395 -0.845 28.725 -0.515 ;
        RECT 28.4 -1.52 28.72 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.755 8.675 30.085 9.005 ;
        RECT 29.755 7.315 30.085 7.645 ;
        RECT 29.755 3.235 30.085 3.565 ;
        RECT 29.755 1.875 30.085 2.205 ;
        RECT 29.755 0.515 30.085 0.845 ;
        RECT 29.755 -0.845 30.085 -0.515 ;
        RECT 29.76 -1.52 30.08 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.115 8.675 31.445 9.005 ;
        RECT 31.115 7.315 31.445 7.645 ;
        RECT 31.115 1.875 31.445 2.205 ;
        RECT 31.115 0.515 31.445 0.845 ;
        RECT 31.115 -0.845 31.445 -0.515 ;
        RECT 31.12 -1.52 31.44 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.475 8.675 32.805 9.005 ;
        RECT 32.475 7.315 32.805 7.645 ;
        RECT 32.475 1.875 32.805 2.205 ;
        RECT 32.475 0.515 32.805 0.845 ;
        RECT 32.475 -0.845 32.805 -0.515 ;
        RECT 32.48 -1.52 32.8 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.835 8.675 34.165 9.005 ;
        RECT 33.835 7.315 34.165 7.645 ;
        RECT 33.835 1.875 34.165 2.205 ;
        RECT 33.835 0.515 34.165 0.845 ;
        RECT 33.835 -0.845 34.165 -0.515 ;
        RECT 33.84 -1.52 34.16 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.195 8.675 35.525 9.005 ;
        RECT 35.195 7.315 35.525 7.645 ;
        RECT 35.195 1.875 35.525 2.205 ;
        RECT 35.195 0.515 35.525 0.845 ;
        RECT 35.195 -0.845 35.525 -0.515 ;
        RECT 35.2 -1.52 35.52 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.555 8.675 36.885 9.005 ;
        RECT 36.555 7.315 36.885 7.645 ;
        RECT 36.555 1.875 36.885 2.205 ;
        RECT 36.555 0.515 36.885 0.845 ;
        RECT 36.555 -0.845 36.885 -0.515 ;
        RECT 36.56 -1.52 36.88 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.915 8.675 38.245 9.005 ;
        RECT 37.915 7.315 38.245 7.645 ;
        RECT 37.915 1.875 38.245 2.205 ;
        RECT 37.915 0.515 38.245 0.845 ;
        RECT 37.915 -0.845 38.245 -0.515 ;
        RECT 37.92 -1.52 38.24 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.275 8.675 39.605 9.005 ;
        RECT 39.275 7.315 39.605 7.645 ;
        RECT 39.275 3.235 39.605 3.565 ;
        RECT 39.275 1.875 39.605 2.205 ;
        RECT 39.275 0.515 39.605 0.845 ;
        RECT 39.275 -0.845 39.605 -0.515 ;
        RECT 39.28 -1.52 39.6 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.635 8.675 40.965 9.005 ;
        RECT 40.635 7.315 40.965 7.645 ;
        RECT 40.635 3.235 40.965 3.565 ;
        RECT 40.635 1.875 40.965 2.205 ;
        RECT 40.635 0.515 40.965 0.845 ;
        RECT 40.635 -0.845 40.965 -0.515 ;
        RECT 40.64 -1.52 40.96 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.995 8.675 42.325 9.005 ;
        RECT 41.995 7.315 42.325 7.645 ;
        RECT 41.995 3.235 42.325 3.565 ;
        RECT 41.995 1.875 42.325 2.205 ;
        RECT 41.995 0.515 42.325 0.845 ;
        RECT 41.995 -0.845 42.325 -0.515 ;
        RECT 42 -1.52 42.32 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.355 8.675 43.685 9.005 ;
        RECT 43.355 7.315 43.685 7.645 ;
        RECT 43.355 1.875 43.685 2.205 ;
        RECT 43.355 0.515 43.685 0.845 ;
        RECT 43.355 -0.845 43.685 -0.515 ;
        RECT 43.36 -1.52 43.68 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.715 8.675 45.045 9.005 ;
        RECT 44.715 7.315 45.045 7.645 ;
        RECT 44.715 1.875 45.045 2.205 ;
        RECT 44.715 0.515 45.045 0.845 ;
        RECT 44.715 -0.845 45.045 -0.515 ;
        RECT 44.72 -1.52 45.04 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.075 8.675 46.405 9.005 ;
        RECT 46.075 7.315 46.405 7.645 ;
        RECT 46.075 1.875 46.405 2.205 ;
        RECT 46.075 0.515 46.405 0.845 ;
        RECT 46.075 -0.845 46.405 -0.515 ;
        RECT 46.08 -1.52 46.4 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.435 8.675 47.765 9.005 ;
        RECT 47.435 7.315 47.765 7.645 ;
        RECT 47.435 1.875 47.765 2.205 ;
        RECT 47.435 0.515 47.765 0.845 ;
        RECT 47.435 -0.845 47.765 -0.515 ;
        RECT 47.44 -1.52 47.76 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.795 8.675 49.125 9.005 ;
        RECT 48.795 7.315 49.125 7.645 ;
        RECT 48.795 1.875 49.125 2.205 ;
        RECT 48.795 0.515 49.125 0.845 ;
        RECT 48.795 -0.845 49.125 -0.515 ;
        RECT 48.8 -1.52 49.12 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.155 8.675 50.485 9.005 ;
        RECT 50.155 7.315 50.485 7.645 ;
        RECT 50.155 1.875 50.485 2.205 ;
        RECT 50.155 0.515 50.485 0.845 ;
        RECT 50.155 -0.845 50.485 -0.515 ;
        RECT 50.16 -1.52 50.48 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.515 8.675 51.845 9.005 ;
        RECT 51.515 7.315 51.845 7.645 ;
        RECT 51.515 3.235 51.845 3.565 ;
        RECT 51.515 1.875 51.845 2.205 ;
        RECT 51.515 0.515 51.845 0.845 ;
        RECT 51.515 -0.845 51.845 -0.515 ;
        RECT 51.52 -1.52 51.84 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.875 8.675 53.205 9.005 ;
        RECT 52.875 7.315 53.205 7.645 ;
        RECT 52.875 3.235 53.205 3.565 ;
        RECT 52.875 1.875 53.205 2.205 ;
        RECT 52.875 0.515 53.205 0.845 ;
        RECT 52.875 -0.845 53.205 -0.515 ;
        RECT 52.88 -1.52 53.2 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.235 8.675 54.565 9.005 ;
        RECT 54.235 7.315 54.565 7.645 ;
        RECT 54.235 3.235 54.565 3.565 ;
        RECT 54.235 1.875 54.565 2.205 ;
        RECT 54.235 0.515 54.565 0.845 ;
        RECT 54.235 -0.845 54.565 -0.515 ;
        RECT 54.24 -1.52 54.56 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.595 8.675 55.925 9.005 ;
        RECT 55.595 7.315 55.925 7.645 ;
        RECT 55.595 1.875 55.925 2.205 ;
        RECT 55.595 0.515 55.925 0.845 ;
        RECT 55.595 -0.845 55.925 -0.515 ;
        RECT 55.6 -1.52 55.92 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.955 8.675 57.285 9.005 ;
        RECT 56.955 7.315 57.285 7.645 ;
        RECT 56.955 1.875 57.285 2.205 ;
        RECT 56.955 0.515 57.285 0.845 ;
        RECT 56.955 -0.845 57.285 -0.515 ;
        RECT 56.96 -1.52 57.28 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.315 8.675 58.645 9.005 ;
        RECT 58.315 7.315 58.645 7.645 ;
        RECT 58.315 1.875 58.645 2.205 ;
        RECT 58.315 0.515 58.645 0.845 ;
        RECT 58.315 -0.845 58.645 -0.515 ;
        RECT 58.32 -1.52 58.64 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.675 8.675 60.005 9.005 ;
        RECT 59.675 7.315 60.005 7.645 ;
        RECT 59.675 1.875 60.005 2.205 ;
        RECT 59.675 0.515 60.005 0.845 ;
        RECT 59.675 -0.845 60.005 -0.515 ;
        RECT 59.68 -1.52 60 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.035 8.675 61.365 9.005 ;
        RECT 61.035 7.315 61.365 7.645 ;
        RECT 61.035 1.875 61.365 2.205 ;
        RECT 61.035 0.515 61.365 0.845 ;
        RECT 61.035 -0.845 61.365 -0.515 ;
        RECT 61.04 -1.52 61.36 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.395 8.675 62.725 9.005 ;
        RECT 62.395 7.315 62.725 7.645 ;
        RECT 62.395 1.875 62.725 2.205 ;
        RECT 62.395 0.515 62.725 0.845 ;
        RECT 62.395 -0.845 62.725 -0.515 ;
        RECT 62.4 -1.52 62.72 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.755 8.675 64.085 9.005 ;
        RECT 63.755 7.315 64.085 7.645 ;
        RECT 63.755 3.235 64.085 3.565 ;
        RECT 63.755 1.875 64.085 2.205 ;
        RECT 63.755 0.515 64.085 0.845 ;
        RECT 63.755 -0.845 64.085 -0.515 ;
        RECT 63.76 -1.52 64.08 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.115 8.675 65.445 9.005 ;
        RECT 65.115 7.315 65.445 7.645 ;
        RECT 65.115 3.235 65.445 3.565 ;
        RECT 65.115 1.875 65.445 2.205 ;
        RECT 65.115 0.515 65.445 0.845 ;
        RECT 65.115 -0.845 65.445 -0.515 ;
        RECT 65.12 -1.52 65.44 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.475 8.675 66.805 9.005 ;
        RECT 66.475 7.315 66.805 7.645 ;
        RECT 66.475 3.235 66.805 3.565 ;
        RECT 66.475 1.875 66.805 2.205 ;
        RECT 66.475 0.515 66.805 0.845 ;
        RECT 66.475 -0.845 66.805 -0.515 ;
        RECT 66.48 -1.52 66.8 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.835 8.675 68.165 9.005 ;
        RECT 67.835 7.315 68.165 7.645 ;
        RECT 67.835 1.875 68.165 2.205 ;
        RECT 67.835 0.515 68.165 0.845 ;
        RECT 67.835 -0.845 68.165 -0.515 ;
        RECT 67.84 -1.52 68.16 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.195 8.675 69.525 9.005 ;
        RECT 69.195 7.315 69.525 7.645 ;
        RECT 69.195 1.875 69.525 2.205 ;
        RECT 69.195 0.515 69.525 0.845 ;
        RECT 69.195 -0.845 69.525 -0.515 ;
        RECT 69.2 -1.52 69.52 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.555 8.675 70.885 9.005 ;
        RECT 70.555 7.315 70.885 7.645 ;
        RECT 70.555 1.875 70.885 2.205 ;
        RECT 70.555 0.515 70.885 0.845 ;
        RECT 70.555 -0.845 70.885 -0.515 ;
        RECT 70.56 -1.52 70.88 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915 8.675 72.245 9.005 ;
        RECT 71.915 7.315 72.245 7.645 ;
        RECT 71.915 1.875 72.245 2.205 ;
        RECT 71.915 0.515 72.245 0.845 ;
        RECT 71.915 -0.845 72.245 -0.515 ;
        RECT 71.92 -1.52 72.24 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.275 8.675 73.605 9.005 ;
        RECT 73.275 7.315 73.605 7.645 ;
        RECT 73.275 1.875 73.605 2.205 ;
        RECT 73.275 0.515 73.605 0.845 ;
        RECT 73.275 -0.845 73.605 -0.515 ;
        RECT 73.28 -1.52 73.6 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.635 8.675 74.965 9.005 ;
        RECT 74.635 7.315 74.965 7.645 ;
        RECT 74.635 1.875 74.965 2.205 ;
        RECT 74.635 0.515 74.965 0.845 ;
        RECT 74.635 -0.845 74.965 -0.515 ;
        RECT 74.64 -1.52 74.96 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.995 8.675 76.325 9.005 ;
        RECT 75.995 7.315 76.325 7.645 ;
        RECT 75.995 3.235 76.325 3.565 ;
        RECT 75.995 1.875 76.325 2.205 ;
        RECT 75.995 0.515 76.325 0.845 ;
        RECT 75.995 -0.845 76.325 -0.515 ;
        RECT 76 -1.52 76.32 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.355 8.675 77.685 9.005 ;
        RECT 77.355 7.315 77.685 7.645 ;
        RECT 77.355 3.235 77.685 3.565 ;
        RECT 77.355 1.875 77.685 2.205 ;
        RECT 77.355 0.515 77.685 0.845 ;
        RECT 77.355 -0.845 77.685 -0.515 ;
        RECT 77.36 -1.52 77.68 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.715 8.675 79.045 9.005 ;
        RECT 78.715 7.315 79.045 7.645 ;
        RECT 78.715 3.235 79.045 3.565 ;
        RECT 78.715 1.875 79.045 2.205 ;
        RECT 78.715 0.515 79.045 0.845 ;
        RECT 78.715 -0.845 79.045 -0.515 ;
        RECT 78.72 -1.52 79.04 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.075 8.675 80.405 9.005 ;
        RECT 80.075 7.315 80.405 7.645 ;
        RECT 80.075 1.875 80.405 2.205 ;
        RECT 80.075 0.515 80.405 0.845 ;
        RECT 80.075 -0.845 80.405 -0.515 ;
        RECT 80.08 -1.52 80.4 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.435 8.675 81.765 9.005 ;
        RECT 81.435 7.315 81.765 7.645 ;
        RECT 81.435 1.875 81.765 2.205 ;
        RECT 81.435 0.515 81.765 0.845 ;
        RECT 81.435 -0.845 81.765 -0.515 ;
        RECT 81.44 -1.52 81.76 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.795 8.675 83.125 9.005 ;
        RECT 82.795 7.315 83.125 7.645 ;
        RECT 82.795 1.875 83.125 2.205 ;
        RECT 82.795 0.515 83.125 0.845 ;
        RECT 82.795 -0.845 83.125 -0.515 ;
        RECT 82.8 -1.52 83.12 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.155 8.675 84.485 9.005 ;
        RECT 84.155 7.315 84.485 7.645 ;
        RECT 84.155 1.875 84.485 2.205 ;
        RECT 84.155 0.515 84.485 0.845 ;
        RECT 84.155 -0.845 84.485 -0.515 ;
        RECT 84.16 -1.52 84.48 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.515 8.675 85.845 9.005 ;
        RECT 85.515 7.315 85.845 7.645 ;
        RECT 85.515 1.875 85.845 2.205 ;
        RECT 85.515 0.515 85.845 0.845 ;
        RECT 85.515 -0.845 85.845 -0.515 ;
        RECT 85.52 -1.52 85.84 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.875 8.675 87.205 9.005 ;
        RECT 86.875 7.315 87.205 7.645 ;
        RECT 86.875 3.235 87.205 3.565 ;
        RECT 86.875 1.875 87.205 2.205 ;
        RECT 86.875 0.515 87.205 0.845 ;
        RECT 86.875 -0.845 87.205 -0.515 ;
        RECT 86.88 -1.52 87.2 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.235 8.675 88.565 9.005 ;
        RECT 88.235 7.315 88.565 7.645 ;
        RECT 88.235 3.235 88.565 3.565 ;
        RECT 88.235 1.875 88.565 2.205 ;
        RECT 88.235 0.515 88.565 0.845 ;
        RECT 88.235 -0.845 88.565 -0.515 ;
        RECT 88.24 -1.52 88.56 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 89.595 8.675 89.925 9.005 ;
        RECT 89.595 7.315 89.925 7.645 ;
        RECT 89.595 3.235 89.925 3.565 ;
        RECT 89.595 1.875 89.925 2.205 ;
        RECT 89.595 0.515 89.925 0.845 ;
        RECT 89.595 -0.845 89.925 -0.515 ;
        RECT 89.6 -1.52 89.92 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.955 8.675 91.285 9.005 ;
        RECT 90.955 7.315 91.285 7.645 ;
        RECT 90.955 1.875 91.285 2.205 ;
        RECT 90.955 0.515 91.285 0.845 ;
        RECT 90.955 -0.845 91.285 -0.515 ;
        RECT 90.96 -1.52 91.28 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.315 8.675 92.645 9.005 ;
        RECT 92.315 7.315 92.645 7.645 ;
        RECT 92.315 1.875 92.645 2.205 ;
        RECT 92.315 0.515 92.645 0.845 ;
        RECT 92.315 -0.845 92.645 -0.515 ;
        RECT 92.32 -1.52 92.64 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.675 8.675 94.005 9.005 ;
        RECT 93.675 7.315 94.005 7.645 ;
        RECT 93.675 1.875 94.005 2.205 ;
        RECT 93.675 0.515 94.005 0.845 ;
        RECT 93.675 -0.845 94.005 -0.515 ;
        RECT 93.68 -1.52 94 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.035 8.675 95.365 9.005 ;
        RECT 95.035 7.315 95.365 7.645 ;
        RECT 95.035 1.875 95.365 2.205 ;
        RECT 95.035 0.515 95.365 0.845 ;
        RECT 95.035 -0.845 95.365 -0.515 ;
        RECT 95.04 -1.52 95.36 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.395 8.675 96.725 9.005 ;
        RECT 96.395 7.315 96.725 7.645 ;
        RECT 96.395 1.875 96.725 2.205 ;
        RECT 96.395 0.515 96.725 0.845 ;
        RECT 96.395 -0.845 96.725 -0.515 ;
        RECT 96.4 -1.52 96.72 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.755 8.675 98.085 9.005 ;
        RECT 97.755 7.315 98.085 7.645 ;
        RECT 97.755 1.875 98.085 2.205 ;
        RECT 97.755 0.515 98.085 0.845 ;
        RECT 97.755 -0.845 98.085 -0.515 ;
        RECT 97.76 -1.52 98.08 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.115 8.675 99.445 9.005 ;
        RECT 99.115 7.315 99.445 7.645 ;
        RECT 99.115 3.235 99.445 3.565 ;
        RECT 99.115 1.875 99.445 2.205 ;
        RECT 99.115 0.515 99.445 0.845 ;
        RECT 99.115 -0.845 99.445 -0.515 ;
        RECT 99.12 -1.52 99.44 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.475 8.675 100.805 9.005 ;
        RECT 100.475 7.315 100.805 7.645 ;
        RECT 100.475 3.235 100.805 3.565 ;
        RECT 100.475 1.875 100.805 2.205 ;
        RECT 100.475 0.515 100.805 0.845 ;
        RECT 100.475 -0.845 100.805 -0.515 ;
        RECT 100.48 -1.52 100.8 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.835 8.675 102.165 9.005 ;
        RECT 101.835 7.315 102.165 7.645 ;
        RECT 101.835 3.235 102.165 3.565 ;
        RECT 101.835 1.875 102.165 2.205 ;
        RECT 101.835 0.515 102.165 0.845 ;
        RECT 101.835 -0.845 102.165 -0.515 ;
        RECT 101.84 -1.52 102.16 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.195 8.675 103.525 9.005 ;
        RECT 103.195 7.315 103.525 7.645 ;
        RECT 103.195 1.875 103.525 2.205 ;
        RECT 103.195 0.515 103.525 0.845 ;
        RECT 103.195 -0.845 103.525 -0.515 ;
        RECT 103.2 -1.52 103.52 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 104.555 8.675 104.885 9.005 ;
        RECT 104.555 7.315 104.885 7.645 ;
        RECT 104.555 1.875 104.885 2.205 ;
        RECT 104.555 0.515 104.885 0.845 ;
        RECT 104.555 -0.845 104.885 -0.515 ;
        RECT 104.56 -1.52 104.88 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.915 8.675 106.245 9.005 ;
        RECT 105.915 7.315 106.245 7.645 ;
        RECT 105.915 1.875 106.245 2.205 ;
        RECT 105.915 0.515 106.245 0.845 ;
        RECT 105.915 -0.845 106.245 -0.515 ;
        RECT 105.92 -1.52 106.24 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.275 8.675 107.605 9.005 ;
        RECT 107.275 7.315 107.605 7.645 ;
        RECT 107.275 1.875 107.605 2.205 ;
        RECT 107.275 0.515 107.605 0.845 ;
        RECT 107.275 -0.845 107.605 -0.515 ;
        RECT 107.28 -1.52 107.6 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.635 8.675 108.965 9.005 ;
        RECT 108.635 7.315 108.965 7.645 ;
        RECT 108.635 1.875 108.965 2.205 ;
        RECT 108.635 0.515 108.965 0.845 ;
        RECT 108.635 -0.845 108.965 -0.515 ;
        RECT 108.64 -1.52 108.96 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.995 8.675 110.325 9.005 ;
        RECT 109.995 7.315 110.325 7.645 ;
        RECT 109.995 1.875 110.325 2.205 ;
        RECT 109.995 0.515 110.325 0.845 ;
        RECT 109.995 -0.845 110.325 -0.515 ;
        RECT 110 -1.52 110.32 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.355 8.675 111.685 9.005 ;
        RECT 111.355 7.315 111.685 7.645 ;
        RECT 111.355 3.235 111.685 3.565 ;
        RECT 111.355 1.875 111.685 2.205 ;
        RECT 111.355 0.515 111.685 0.845 ;
        RECT 111.355 -0.845 111.685 -0.515 ;
        RECT 111.36 -1.52 111.68 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.715 8.675 113.045 9.005 ;
        RECT 112.715 7.315 113.045 7.645 ;
        RECT 112.715 3.235 113.045 3.565 ;
        RECT 112.715 1.875 113.045 2.205 ;
        RECT 112.715 0.515 113.045 0.845 ;
        RECT 112.715 -0.845 113.045 -0.515 ;
        RECT 112.72 -1.52 113.04 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.075 8.675 114.405 9.005 ;
        RECT 114.075 7.315 114.405 7.645 ;
        RECT 114.075 3.235 114.405 3.565 ;
        RECT 114.075 1.875 114.405 2.205 ;
        RECT 114.075 0.515 114.405 0.845 ;
        RECT 114.075 -0.845 114.405 -0.515 ;
        RECT 114.08 -1.52 114.4 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.435 8.675 115.765 9.005 ;
        RECT 115.435 7.315 115.765 7.645 ;
        RECT 115.435 1.875 115.765 2.205 ;
        RECT 115.435 0.515 115.765 0.845 ;
        RECT 115.435 -0.845 115.765 -0.515 ;
        RECT 115.44 -1.52 115.76 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.795 8.675 117.125 9.005 ;
        RECT 116.795 7.315 117.125 7.645 ;
        RECT 116.795 1.875 117.125 2.205 ;
        RECT 116.795 0.515 117.125 0.845 ;
        RECT 116.795 -0.845 117.125 -0.515 ;
        RECT 116.8 -1.52 117.12 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.155 8.675 118.485 9.005 ;
        RECT 118.155 7.315 118.485 7.645 ;
        RECT 118.155 1.875 118.485 2.205 ;
        RECT 118.155 0.515 118.485 0.845 ;
        RECT 118.155 -0.845 118.485 -0.515 ;
        RECT 118.16 -1.52 118.48 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 119.515 8.675 119.845 9.005 ;
        RECT 119.515 7.315 119.845 7.645 ;
        RECT 119.515 1.875 119.845 2.205 ;
        RECT 119.515 0.515 119.845 0.845 ;
        RECT 119.515 -0.845 119.845 -0.515 ;
        RECT 119.52 -1.52 119.84 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.875 8.675 121.205 9.005 ;
        RECT 120.875 7.315 121.205 7.645 ;
        RECT 120.875 1.875 121.205 2.205 ;
        RECT 120.875 0.515 121.205 0.845 ;
        RECT 120.875 -0.845 121.205 -0.515 ;
        RECT 120.88 -1.52 121.2 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.235 8.675 122.565 9.005 ;
        RECT 122.235 7.315 122.565 7.645 ;
        RECT 122.235 1.875 122.565 2.205 ;
        RECT 122.235 0.515 122.565 0.845 ;
        RECT 122.235 -0.845 122.565 -0.515 ;
        RECT 122.24 -1.52 122.56 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.595 8.675 123.925 9.005 ;
        RECT 123.595 7.315 123.925 7.645 ;
        RECT 123.595 3.235 123.925 3.565 ;
        RECT 123.595 1.875 123.925 2.205 ;
        RECT 123.595 0.515 123.925 0.845 ;
        RECT 123.595 -0.845 123.925 -0.515 ;
        RECT 123.6 -1.52 123.92 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.955 8.675 125.285 9.005 ;
        RECT 124.955 7.315 125.285 7.645 ;
        RECT 124.955 3.235 125.285 3.565 ;
        RECT 124.955 1.875 125.285 2.205 ;
        RECT 124.955 0.515 125.285 0.845 ;
        RECT 124.955 -0.845 125.285 -0.515 ;
        RECT 124.96 -1.52 125.28 9.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.315 0.515 126.645 0.845 ;
        RECT 126.315 -0.845 126.645 -0.515 ;
        RECT 126.32 -1.52 126.64 9.005 ;
        RECT 126.315 8.675 126.645 9.005 ;
        RECT 126.315 7.315 126.645 7.645 ;
        RECT 126.315 3.235 126.645 3.565 ;
        RECT 126.315 1.875 126.645 2.205 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 547.235 7.995 547.565 8.325 ;
        RECT 547.235 2.555 547.565 2.885 ;
        RECT 547.235 1.195 547.565 1.525 ;
        RECT 547.235 -0.165 547.565 0.165 ;
        RECT 547.235 -1.525 547.565 -1.195 ;
        RECT 547.24 -1.525 547.56 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 548.595 7.995 548.925 8.325 ;
        RECT 548.595 2.555 548.925 2.885 ;
        RECT 548.595 1.195 548.925 1.525 ;
        RECT 548.595 -0.165 548.925 0.165 ;
        RECT 548.595 -1.525 548.925 -1.195 ;
        RECT 548.6 -1.525 548.92 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 549.955 7.995 550.285 8.325 ;
        RECT 549.955 2.555 550.285 2.885 ;
        RECT 549.955 1.195 550.285 1.525 ;
        RECT 549.955 -0.165 550.285 0.165 ;
        RECT 549.955 -1.525 550.285 -1.195 ;
        RECT 549.96 -1.525 550.28 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 551.315 7.995 551.645 8.325 ;
        RECT 551.315 2.555 551.645 2.885 ;
        RECT 551.315 1.195 551.645 1.525 ;
        RECT 551.315 -0.165 551.645 0.165 ;
        RECT 551.315 -1.525 551.645 -1.195 ;
        RECT 551.32 -1.525 551.64 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 552.675 7.995 553.005 8.325 ;
        RECT 552.675 2.555 553.005 2.885 ;
        RECT 552.675 1.195 553.005 1.525 ;
        RECT 552.675 -0.165 553.005 0.165 ;
        RECT 552.675 -1.525 553.005 -1.195 ;
        RECT 552.68 -1.525 553 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 554.035 7.995 554.365 8.325 ;
        RECT 554.035 2.555 554.365 2.885 ;
        RECT 554.035 1.195 554.365 1.525 ;
        RECT 554.035 -0.165 554.365 0.165 ;
        RECT 554.035 -1.525 554.365 -1.195 ;
        RECT 554.04 -1.525 554.36 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 555.395 7.995 555.725 8.325 ;
        RECT 555.395 2.555 555.725 2.885 ;
        RECT 555.395 1.195 555.725 1.525 ;
        RECT 555.395 -0.165 555.725 0.165 ;
        RECT 555.395 -1.525 555.725 -1.195 ;
        RECT 555.4 -1.525 555.72 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 556.755 7.995 557.085 8.325 ;
        RECT 556.755 2.555 557.085 2.885 ;
        RECT 556.755 1.195 557.085 1.525 ;
        RECT 556.755 -0.165 557.085 0.165 ;
        RECT 556.755 -1.525 557.085 -1.195 ;
        RECT 556.76 -1.525 557.08 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 558.115 7.995 558.445 8.325 ;
        RECT 558.115 2.555 558.445 2.885 ;
        RECT 558.115 1.195 558.445 1.525 ;
        RECT 558.115 -0.165 558.445 0.165 ;
        RECT 558.115 -1.525 558.445 -1.195 ;
        RECT 558.12 -1.525 558.44 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 559.475 7.995 559.805 8.325 ;
        RECT 559.475 2.555 559.805 2.885 ;
        RECT 559.475 1.195 559.805 1.525 ;
        RECT 559.475 -0.165 559.805 0.165 ;
        RECT 559.475 -1.525 559.805 -1.195 ;
        RECT 559.48 -1.525 559.8 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 560.835 7.995 561.165 8.325 ;
        RECT 560.835 2.555 561.165 2.885 ;
        RECT 560.835 1.195 561.165 1.525 ;
        RECT 560.835 -0.165 561.165 0.165 ;
        RECT 560.835 -1.525 561.165 -1.195 ;
        RECT 560.84 -1.525 561.16 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 562.195 7.995 562.525 8.325 ;
        RECT 562.195 2.555 562.525 2.885 ;
        RECT 562.195 1.195 562.525 1.525 ;
        RECT 562.195 -0.165 562.525 0.165 ;
        RECT 562.195 -1.525 562.525 -1.195 ;
        RECT 562.2 -1.525 562.52 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 563.555 7.995 563.885 8.325 ;
        RECT 563.555 2.555 563.885 2.885 ;
        RECT 563.555 1.195 563.885 1.525 ;
        RECT 563.555 -0.165 563.885 0.165 ;
        RECT 563.555 -1.525 563.885 -1.195 ;
        RECT 563.56 -1.525 563.88 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 564.915 7.995 565.245 8.325 ;
        RECT 564.915 2.555 565.245 2.885 ;
        RECT 564.915 1.195 565.245 1.525 ;
        RECT 564.915 -0.165 565.245 0.165 ;
        RECT 564.915 -1.525 565.245 -1.195 ;
        RECT 564.92 -1.525 565.24 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 566.275 7.995 566.605 8.325 ;
        RECT 566.275 2.555 566.605 2.885 ;
        RECT 566.275 1.195 566.605 1.525 ;
        RECT 566.275 -0.165 566.605 0.165 ;
        RECT 566.275 -1.525 566.605 -1.195 ;
        RECT 566.28 -1.525 566.6 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 567.635 7.995 567.965 8.325 ;
        RECT 567.635 2.555 567.965 2.885 ;
        RECT 567.635 1.195 567.965 1.525 ;
        RECT 567.635 -0.165 567.965 0.165 ;
        RECT 567.635 -1.525 567.965 -1.195 ;
        RECT 567.64 -1.525 567.96 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 568.995 7.995 569.325 8.325 ;
        RECT 568.995 2.555 569.325 2.885 ;
        RECT 568.995 1.195 569.325 1.525 ;
        RECT 568.995 -0.165 569.325 0.165 ;
        RECT 568.995 -1.525 569.325 -1.195 ;
        RECT 569 -1.525 569.32 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 570.355 7.995 570.685 8.325 ;
        RECT 570.355 2.555 570.685 2.885 ;
        RECT 570.355 1.195 570.685 1.525 ;
        RECT 570.355 -0.165 570.685 0.165 ;
        RECT 570.355 -1.525 570.685 -1.195 ;
        RECT 570.36 -1.525 570.68 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 571.715 7.995 572.045 8.325 ;
        RECT 571.715 2.555 572.045 2.885 ;
        RECT 571.715 1.195 572.045 1.525 ;
        RECT 571.715 -0.165 572.045 0.165 ;
        RECT 571.715 -1.525 572.045 -1.195 ;
        RECT 571.72 -1.525 572.04 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 573.075 7.995 573.405 8.325 ;
        RECT 573.075 2.555 573.405 2.885 ;
        RECT 573.075 1.195 573.405 1.525 ;
        RECT 573.075 -0.165 573.405 0.165 ;
        RECT 573.075 -1.525 573.405 -1.195 ;
        RECT 573.08 -1.525 573.4 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 574.435 7.995 574.765 8.325 ;
        RECT 574.435 2.555 574.765 2.885 ;
        RECT 574.435 1.195 574.765 1.525 ;
        RECT 574.435 -0.165 574.765 0.165 ;
        RECT 574.435 -1.525 574.765 -1.195 ;
        RECT 574.44 -1.525 574.76 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 575.795 7.995 576.125 8.325 ;
        RECT 575.795 2.555 576.125 2.885 ;
        RECT 575.795 1.195 576.125 1.525 ;
        RECT 575.795 -0.165 576.125 0.165 ;
        RECT 575.795 -1.525 576.125 -1.195 ;
        RECT 575.8 -1.525 576.12 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 577.155 7.995 577.485 8.325 ;
        RECT 577.155 2.555 577.485 2.885 ;
        RECT 577.155 1.195 577.485 1.525 ;
        RECT 577.155 -0.165 577.485 0.165 ;
        RECT 577.155 -1.525 577.485 -1.195 ;
        RECT 577.16 -1.525 577.48 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 578.515 7.995 578.845 8.325 ;
        RECT 578.515 2.555 578.845 2.885 ;
        RECT 578.515 1.195 578.845 1.525 ;
        RECT 578.515 -0.165 578.845 0.165 ;
        RECT 578.515 -1.525 578.845 -1.195 ;
        RECT 578.52 -1.525 578.84 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 579.875 7.995 580.205 8.325 ;
        RECT 579.875 2.555 580.205 2.885 ;
        RECT 579.875 1.195 580.205 1.525 ;
        RECT 579.875 -0.165 580.205 0.165 ;
        RECT 579.875 -1.525 580.205 -1.195 ;
        RECT 579.88 -1.525 580.2 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 581.235 7.995 581.565 8.325 ;
        RECT 581.235 2.555 581.565 2.885 ;
        RECT 581.235 1.195 581.565 1.525 ;
        RECT 581.235 -0.165 581.565 0.165 ;
        RECT 581.235 -1.525 581.565 -1.195 ;
        RECT 581.24 -1.525 581.56 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 582.595 7.995 582.925 8.325 ;
        RECT 582.595 2.555 582.925 2.885 ;
        RECT 582.595 1.195 582.925 1.525 ;
        RECT 582.595 -0.165 582.925 0.165 ;
        RECT 582.595 -1.525 582.925 -1.195 ;
        RECT 582.6 -1.525 582.92 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 583.955 7.995 584.285 8.325 ;
        RECT 583.955 2.555 584.285 2.885 ;
        RECT 583.955 1.195 584.285 1.525 ;
        RECT 583.955 -0.165 584.285 0.165 ;
        RECT 583.955 -1.525 584.285 -1.195 ;
        RECT 583.96 -1.525 584.28 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 585.315 7.995 585.645 8.325 ;
        RECT 585.315 2.555 585.645 2.885 ;
        RECT 585.315 1.195 585.645 1.525 ;
        RECT 585.315 -0.165 585.645 0.165 ;
        RECT 585.315 -1.525 585.645 -1.195 ;
        RECT 585.32 -1.525 585.64 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 586.675 7.995 587.005 8.325 ;
        RECT 586.675 2.555 587.005 2.885 ;
        RECT 586.675 1.195 587.005 1.525 ;
        RECT 586.675 -0.165 587.005 0.165 ;
        RECT 586.675 -1.525 587.005 -1.195 ;
        RECT 586.68 -1.525 587 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 588.035 7.995 588.365 8.325 ;
        RECT 588.035 2.555 588.365 2.885 ;
        RECT 588.035 1.195 588.365 1.525 ;
        RECT 588.035 -0.165 588.365 0.165 ;
        RECT 588.035 -1.525 588.365 -1.195 ;
        RECT 588.04 -1.525 588.36 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 589.395 7.995 589.725 8.325 ;
        RECT 589.395 2.555 589.725 2.885 ;
        RECT 589.395 1.195 589.725 1.525 ;
        RECT 589.395 -0.165 589.725 0.165 ;
        RECT 589.395 -1.525 589.725 -1.195 ;
        RECT 589.4 -1.525 589.72 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 590.755 7.995 591.085 8.325 ;
        RECT 590.755 2.555 591.085 2.885 ;
        RECT 590.755 1.195 591.085 1.525 ;
        RECT 590.755 -0.165 591.085 0.165 ;
        RECT 590.755 -1.525 591.085 -1.195 ;
        RECT 590.76 -1.525 591.08 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 592.115 7.995 592.445 8.325 ;
        RECT 592.115 2.555 592.445 2.885 ;
        RECT 592.115 1.195 592.445 1.525 ;
        RECT 592.115 -0.165 592.445 0.165 ;
        RECT 592.115 -1.525 592.445 -1.195 ;
        RECT 592.12 -1.525 592.44 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 593.475 7.995 593.805 8.325 ;
        RECT 593.475 2.555 593.805 2.885 ;
        RECT 593.475 1.195 593.805 1.525 ;
        RECT 593.475 -0.165 593.805 0.165 ;
        RECT 593.475 -1.525 593.805 -1.195 ;
        RECT 593.48 -1.525 593.8 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 594.835 7.995 595.165 8.325 ;
        RECT 594.835 2.555 595.165 2.885 ;
        RECT 594.835 1.195 595.165 1.525 ;
        RECT 594.835 -0.165 595.165 0.165 ;
        RECT 594.835 -1.525 595.165 -1.195 ;
        RECT 594.84 -1.525 595.16 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 596.195 7.995 596.525 8.325 ;
        RECT 596.195 2.555 596.525 2.885 ;
        RECT 596.195 1.195 596.525 1.525 ;
        RECT 596.195 -0.165 596.525 0.165 ;
        RECT 596.195 -1.525 596.525 -1.195 ;
        RECT 596.2 -1.525 596.52 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 597.555 7.995 597.885 8.325 ;
        RECT 597.555 2.555 597.885 2.885 ;
        RECT 597.555 1.195 597.885 1.525 ;
        RECT 597.555 -0.165 597.885 0.165 ;
        RECT 597.555 -1.525 597.885 -1.195 ;
        RECT 597.56 -1.525 597.88 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 598.915 7.995 599.245 8.325 ;
        RECT 598.915 2.555 599.245 2.885 ;
        RECT 598.915 1.195 599.245 1.525 ;
        RECT 598.915 -0.165 599.245 0.165 ;
        RECT 598.915 -1.525 599.245 -1.195 ;
        RECT 598.92 -1.525 599.24 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 600.275 7.995 600.605 8.325 ;
        RECT 600.275 2.555 600.605 2.885 ;
        RECT 600.275 1.195 600.605 1.525 ;
        RECT 600.275 -0.165 600.605 0.165 ;
        RECT 600.275 -1.525 600.605 -1.195 ;
        RECT 600.28 -1.525 600.6 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 601.635 7.995 601.965 8.325 ;
        RECT 601.635 2.555 601.965 2.885 ;
        RECT 601.635 1.195 601.965 1.525 ;
        RECT 601.635 -0.165 601.965 0.165 ;
        RECT 601.635 -1.525 601.965 -1.195 ;
        RECT 601.64 -1.525 601.96 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 602.995 7.995 603.325 8.325 ;
        RECT 602.995 2.555 603.325 2.885 ;
        RECT 602.995 1.195 603.325 1.525 ;
        RECT 602.995 -0.165 603.325 0.165 ;
        RECT 602.995 -1.525 603.325 -1.195 ;
        RECT 603 -1.525 603.32 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 604.355 7.995 604.685 8.325 ;
        RECT 604.355 2.555 604.685 2.885 ;
        RECT 604.355 1.195 604.685 1.525 ;
        RECT 604.355 -0.165 604.685 0.165 ;
        RECT 604.355 -1.525 604.685 -1.195 ;
        RECT 604.36 -1.525 604.68 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 605.715 7.995 606.045 8.325 ;
        RECT 605.715 2.555 606.045 2.885 ;
        RECT 605.715 1.195 606.045 1.525 ;
        RECT 605.715 -0.165 606.045 0.165 ;
        RECT 605.715 -1.525 606.045 -1.195 ;
        RECT 605.72 -1.525 606.04 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 607.075 7.995 607.405 8.325 ;
        RECT 607.075 2.555 607.405 2.885 ;
        RECT 607.075 1.195 607.405 1.525 ;
        RECT 607.075 -0.165 607.405 0.165 ;
        RECT 607.075 -1.525 607.405 -1.195 ;
        RECT 607.08 -1.525 607.4 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 608.435 7.995 608.765 8.325 ;
        RECT 608.435 2.555 608.765 2.885 ;
        RECT 608.435 1.195 608.765 1.525 ;
        RECT 608.435 -0.165 608.765 0.165 ;
        RECT 608.435 -1.525 608.765 -1.195 ;
        RECT 608.44 -1.525 608.76 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 609.795 7.995 610.125 8.325 ;
        RECT 609.795 2.555 610.125 2.885 ;
        RECT 609.795 1.195 610.125 1.525 ;
        RECT 609.795 -0.165 610.125 0.165 ;
        RECT 609.795 -1.525 610.125 -1.195 ;
        RECT 609.8 -1.525 610.12 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 611.155 7.995 611.485 8.325 ;
        RECT 611.155 2.555 611.485 2.885 ;
        RECT 611.155 1.195 611.485 1.525 ;
        RECT 611.155 -0.165 611.485 0.165 ;
        RECT 611.155 -1.525 611.485 -1.195 ;
        RECT 611.16 -1.525 611.48 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 612.515 7.995 612.845 8.325 ;
        RECT 612.515 2.555 612.845 2.885 ;
        RECT 612.515 1.195 612.845 1.525 ;
        RECT 612.515 -0.165 612.845 0.165 ;
        RECT 612.515 -1.525 612.845 -1.195 ;
        RECT 612.52 -1.525 612.84 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 613.875 7.995 614.205 8.325 ;
        RECT 613.875 2.555 614.205 2.885 ;
        RECT 613.875 1.195 614.205 1.525 ;
        RECT 613.875 -0.165 614.205 0.165 ;
        RECT 613.875 -1.525 614.205 -1.195 ;
        RECT 613.88 -1.525 614.2 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 615.235 7.995 615.565 8.325 ;
        RECT 615.235 2.555 615.565 2.885 ;
        RECT 615.235 1.195 615.565 1.525 ;
        RECT 615.235 -0.165 615.565 0.165 ;
        RECT 615.235 -1.525 615.565 -1.195 ;
        RECT 615.24 -1.525 615.56 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 616.595 7.995 616.925 8.325 ;
        RECT 616.595 2.555 616.925 2.885 ;
        RECT 616.595 1.195 616.925 1.525 ;
        RECT 616.595 -0.165 616.925 0.165 ;
        RECT 616.595 -1.525 616.925 -1.195 ;
        RECT 616.6 -1.525 616.92 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 617.955 7.995 618.285 8.325 ;
        RECT 617.955 2.555 618.285 2.885 ;
        RECT 617.955 1.195 618.285 1.525 ;
        RECT 617.955 -0.165 618.285 0.165 ;
        RECT 617.955 -1.525 618.285 -1.195 ;
        RECT 617.96 -1.525 618.28 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 619.315 7.995 619.645 8.325 ;
        RECT 619.315 2.555 619.645 2.885 ;
        RECT 619.315 1.195 619.645 1.525 ;
        RECT 619.315 -0.165 619.645 0.165 ;
        RECT 619.315 -1.525 619.645 -1.195 ;
        RECT 619.32 -1.525 619.64 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 620.675 7.995 621.005 8.325 ;
        RECT 620.675 2.555 621.005 2.885 ;
        RECT 620.675 1.195 621.005 1.525 ;
        RECT 620.675 -0.165 621.005 0.165 ;
        RECT 620.675 -1.525 621.005 -1.195 ;
        RECT 620.68 -1.525 621 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 622.035 7.995 622.365 8.325 ;
        RECT 622.035 2.555 622.365 2.885 ;
        RECT 622.035 1.195 622.365 1.525 ;
        RECT 622.035 -0.165 622.365 0.165 ;
        RECT 622.035 -1.525 622.365 -1.195 ;
        RECT 622.04 -1.525 622.36 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 623.395 7.995 623.725 8.325 ;
        RECT 623.395 2.555 623.725 2.885 ;
        RECT 623.395 1.195 623.725 1.525 ;
        RECT 623.395 -0.165 623.725 0.165 ;
        RECT 623.395 -1.525 623.725 -1.195 ;
        RECT 623.4 -1.525 623.72 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 624.755 7.995 625.085 8.325 ;
        RECT 624.755 2.555 625.085 2.885 ;
        RECT 624.755 1.195 625.085 1.525 ;
        RECT 624.755 -0.165 625.085 0.165 ;
        RECT 624.755 -1.525 625.085 -1.195 ;
        RECT 624.76 -1.525 625.08 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 626.115 7.995 626.445 8.325 ;
        RECT 626.115 2.555 626.445 2.885 ;
        RECT 626.115 1.195 626.445 1.525 ;
        RECT 626.115 -0.165 626.445 0.165 ;
        RECT 626.115 -1.525 626.445 -1.195 ;
        RECT 626.12 -1.525 626.44 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 627.475 7.995 627.805 8.325 ;
        RECT 627.475 2.555 627.805 2.885 ;
        RECT 627.475 1.195 627.805 1.525 ;
        RECT 627.475 -0.165 627.805 0.165 ;
        RECT 627.475 -1.525 627.805 -1.195 ;
        RECT 627.48 -1.525 627.8 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 628.835 7.995 629.165 8.325 ;
        RECT 628.835 2.555 629.165 2.885 ;
        RECT 628.835 1.195 629.165 1.525 ;
        RECT 628.835 -0.165 629.165 0.165 ;
        RECT 628.835 -1.525 629.165 -1.195 ;
        RECT 628.84 -1.525 629.16 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 630.195 7.995 630.525 8.325 ;
        RECT 630.195 2.555 630.525 2.885 ;
        RECT 630.195 1.195 630.525 1.525 ;
        RECT 630.195 -0.165 630.525 0.165 ;
        RECT 630.195 -1.525 630.525 -1.195 ;
        RECT 630.2 -1.525 630.52 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 631.555 7.995 631.885 8.325 ;
        RECT 631.555 2.555 631.885 2.885 ;
        RECT 631.555 1.195 631.885 1.525 ;
        RECT 631.555 -0.165 631.885 0.165 ;
        RECT 631.555 -1.525 631.885 -1.195 ;
        RECT 631.56 -1.525 631.88 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 632.915 7.995 633.245 8.325 ;
        RECT 632.915 2.555 633.245 2.885 ;
        RECT 632.915 1.195 633.245 1.525 ;
        RECT 632.915 -0.165 633.245 0.165 ;
        RECT 632.915 -1.525 633.245 -1.195 ;
        RECT 632.92 -1.525 633.24 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 634.275 7.995 634.605 8.325 ;
        RECT 634.275 2.555 634.605 2.885 ;
        RECT 634.275 1.195 634.605 1.525 ;
        RECT 634.275 -0.165 634.605 0.165 ;
        RECT 634.275 -1.525 634.605 -1.195 ;
        RECT 634.28 -1.525 634.6 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 635.635 7.995 635.965 8.325 ;
        RECT 635.635 2.555 635.965 2.885 ;
        RECT 635.635 1.195 635.965 1.525 ;
        RECT 635.635 -0.165 635.965 0.165 ;
        RECT 635.635 -1.525 635.965 -1.195 ;
        RECT 635.64 -1.525 635.96 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 636.995 7.995 637.325 8.325 ;
        RECT 636.995 2.555 637.325 2.885 ;
        RECT 636.995 1.195 637.325 1.525 ;
        RECT 636.995 -0.165 637.325 0.165 ;
        RECT 636.995 -1.525 637.325 -1.195 ;
        RECT 637 -1.525 637.32 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 638.355 7.995 638.685 8.325 ;
        RECT 638.355 2.555 638.685 2.885 ;
        RECT 638.355 1.195 638.685 1.525 ;
        RECT 638.355 -0.165 638.685 0.165 ;
        RECT 638.355 -1.525 638.685 -1.195 ;
        RECT 638.36 -1.525 638.68 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 639.715 7.995 640.045 8.325 ;
        RECT 639.715 2.555 640.045 2.885 ;
        RECT 639.715 1.195 640.045 1.525 ;
        RECT 639.715 -0.165 640.045 0.165 ;
        RECT 639.715 -1.525 640.045 -1.195 ;
        RECT 639.72 -1.525 640.04 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 641.075 7.995 641.405 8.325 ;
        RECT 641.075 2.555 641.405 2.885 ;
        RECT 641.075 1.195 641.405 1.525 ;
        RECT 641.075 -0.165 641.405 0.165 ;
        RECT 641.075 -1.525 641.405 -1.195 ;
        RECT 641.08 -1.525 641.4 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 642.435 7.995 642.765 8.325 ;
        RECT 642.435 2.555 642.765 2.885 ;
        RECT 642.435 1.195 642.765 1.525 ;
        RECT 642.435 -0.165 642.765 0.165 ;
        RECT 642.435 -1.525 642.765 -1.195 ;
        RECT 642.44 -1.525 642.76 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 643.795 7.995 644.125 8.325 ;
        RECT 643.795 2.555 644.125 2.885 ;
        RECT 643.795 1.195 644.125 1.525 ;
        RECT 643.795 -0.165 644.125 0.165 ;
        RECT 643.795 -1.525 644.125 -1.195 ;
        RECT 643.8 -1.525 644.12 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 645.155 7.995 645.485 8.325 ;
        RECT 645.155 2.555 645.485 2.885 ;
        RECT 645.155 1.195 645.485 1.525 ;
        RECT 645.155 -0.165 645.485 0.165 ;
        RECT 645.155 -1.525 645.485 -1.195 ;
        RECT 645.16 -1.525 645.48 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 646.515 7.995 646.845 8.325 ;
        RECT 646.515 2.555 646.845 2.885 ;
        RECT 646.515 1.195 646.845 1.525 ;
        RECT 646.515 -0.165 646.845 0.165 ;
        RECT 646.515 -1.525 646.845 -1.195 ;
        RECT 646.52 -1.525 646.84 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 647.875 7.995 648.205 8.325 ;
        RECT 647.875 2.555 648.205 2.885 ;
        RECT 647.875 1.195 648.205 1.525 ;
        RECT 647.875 -0.165 648.205 0.165 ;
        RECT 647.875 -1.525 648.205 -1.195 ;
        RECT 647.88 -1.525 648.2 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 649.235 7.995 649.565 8.325 ;
        RECT 649.235 2.555 649.565 2.885 ;
        RECT 649.235 1.195 649.565 1.525 ;
        RECT 649.235 -0.165 649.565 0.165 ;
        RECT 649.235 -1.525 649.565 -1.195 ;
        RECT 649.24 -1.525 649.56 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 650.595 7.995 650.925 8.325 ;
        RECT 650.595 2.555 650.925 2.885 ;
        RECT 650.595 1.195 650.925 1.525 ;
        RECT 650.595 -0.165 650.925 0.165 ;
        RECT 650.595 -1.525 650.925 -1.195 ;
        RECT 650.6 -1.525 650.92 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 651.955 7.995 652.285 8.325 ;
        RECT 651.955 2.555 652.285 2.885 ;
        RECT 651.955 1.195 652.285 1.525 ;
        RECT 651.955 -0.165 652.285 0.165 ;
        RECT 651.955 -1.525 652.285 -1.195 ;
        RECT 651.96 -1.525 652.28 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 653.315 7.995 653.645 8.325 ;
        RECT 653.315 2.555 653.645 2.885 ;
        RECT 653.315 1.195 653.645 1.525 ;
        RECT 653.315 -0.165 653.645 0.165 ;
        RECT 653.315 -1.525 653.645 -1.195 ;
        RECT 653.32 -1.525 653.64 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 654.675 7.995 655.005 8.325 ;
        RECT 654.675 2.555 655.005 2.885 ;
        RECT 654.675 1.195 655.005 1.525 ;
        RECT 654.675 -0.165 655.005 0.165 ;
        RECT 654.675 -1.525 655.005 -1.195 ;
        RECT 654.68 -1.525 655 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 656.035 7.995 656.365 8.325 ;
        RECT 656.035 2.555 656.365 2.885 ;
        RECT 656.035 1.195 656.365 1.525 ;
        RECT 656.035 -0.165 656.365 0.165 ;
        RECT 656.035 -1.525 656.365 -1.195 ;
        RECT 656.04 -1.525 656.36 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 657.395 7.995 657.725 8.325 ;
        RECT 657.395 2.555 657.725 2.885 ;
        RECT 657.395 1.195 657.725 1.525 ;
        RECT 657.395 -0.165 657.725 0.165 ;
        RECT 657.395 -1.525 657.725 -1.195 ;
        RECT 657.4 -1.525 657.72 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 658.755 7.995 659.085 8.325 ;
        RECT 658.755 2.555 659.085 2.885 ;
        RECT 658.755 1.195 659.085 1.525 ;
        RECT 658.755 -0.165 659.085 0.165 ;
        RECT 658.755 -1.525 659.085 -1.195 ;
        RECT 658.76 -1.525 659.08 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 660.115 7.995 660.445 8.325 ;
        RECT 660.115 2.555 660.445 2.885 ;
        RECT 660.115 1.195 660.445 1.525 ;
        RECT 660.115 -0.165 660.445 0.165 ;
        RECT 660.115 -1.525 660.445 -1.195 ;
        RECT 660.12 -1.525 660.44 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 661.475 7.995 661.805 8.325 ;
        RECT 661.475 2.555 661.805 2.885 ;
        RECT 661.475 1.195 661.805 1.525 ;
        RECT 661.475 -0.165 661.805 0.165 ;
        RECT 661.475 -1.525 661.805 -1.195 ;
        RECT 661.48 -1.525 661.8 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 662.835 7.995 663.165 8.325 ;
        RECT 662.835 2.555 663.165 2.885 ;
        RECT 662.835 1.195 663.165 1.525 ;
        RECT 662.835 -0.165 663.165 0.165 ;
        RECT 662.835 -1.525 663.165 -1.195 ;
        RECT 662.84 -1.525 663.16 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 664.195 7.995 664.525 8.325 ;
        RECT 664.195 2.555 664.525 2.885 ;
        RECT 664.195 1.195 664.525 1.525 ;
        RECT 664.195 -0.165 664.525 0.165 ;
        RECT 664.195 -1.525 664.525 -1.195 ;
        RECT 664.2 -1.525 664.52 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 665.555 7.995 665.885 8.325 ;
        RECT 665.555 2.555 665.885 2.885 ;
        RECT 665.555 1.195 665.885 1.525 ;
        RECT 665.555 -0.165 665.885 0.165 ;
        RECT 665.555 -1.525 665.885 -1.195 ;
        RECT 665.56 -1.525 665.88 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 666.915 7.995 667.245 8.325 ;
        RECT 666.915 2.555 667.245 2.885 ;
        RECT 666.915 1.195 667.245 1.525 ;
        RECT 666.915 -0.165 667.245 0.165 ;
        RECT 666.915 -1.525 667.245 -1.195 ;
        RECT 666.92 -1.525 667.24 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 668.275 7.995 668.605 8.325 ;
        RECT 668.275 2.555 668.605 2.885 ;
        RECT 668.275 1.195 668.605 1.525 ;
        RECT 668.275 -0.165 668.605 0.165 ;
        RECT 668.275 -1.525 668.605 -1.195 ;
        RECT 668.28 -1.525 668.6 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 669.635 7.995 669.965 8.325 ;
        RECT 669.635 2.555 669.965 2.885 ;
        RECT 669.635 1.195 669.965 1.525 ;
        RECT 669.635 -0.165 669.965 0.165 ;
        RECT 669.635 -1.525 669.965 -1.195 ;
        RECT 669.64 -1.525 669.96 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 670.995 7.995 671.325 8.325 ;
        RECT 670.995 2.555 671.325 2.885 ;
        RECT 670.995 1.195 671.325 1.525 ;
        RECT 670.995 -0.165 671.325 0.165 ;
        RECT 670.995 -1.525 671.325 -1.195 ;
        RECT 671 -1.525 671.32 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 672.355 7.995 672.685 8.325 ;
        RECT 672.355 2.555 672.685 2.885 ;
        RECT 672.355 1.195 672.685 1.525 ;
        RECT 672.355 -0.165 672.685 0.165 ;
        RECT 672.355 -1.525 672.685 -1.195 ;
        RECT 672.36 -1.525 672.68 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 673.715 7.995 674.045 8.325 ;
        RECT 673.715 2.555 674.045 2.885 ;
        RECT 673.715 1.195 674.045 1.525 ;
        RECT 673.715 -0.165 674.045 0.165 ;
        RECT 673.715 -1.525 674.045 -1.195 ;
        RECT 673.72 -1.525 674.04 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 675.075 7.995 675.405 8.325 ;
        RECT 675.075 2.555 675.405 2.885 ;
        RECT 675.075 1.195 675.405 1.525 ;
        RECT 675.075 -0.165 675.405 0.165 ;
        RECT 675.075 -1.525 675.405 -1.195 ;
        RECT 675.08 -1.525 675.4 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 676.435 7.995 676.765 8.325 ;
        RECT 676.435 2.555 676.765 2.885 ;
        RECT 676.435 1.195 676.765 1.525 ;
        RECT 676.435 -0.165 676.765 0.165 ;
        RECT 676.435 -1.525 676.765 -1.195 ;
        RECT 676.44 -1.525 676.76 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 677.795 7.995 678.125 8.325 ;
        RECT 677.795 2.555 678.125 2.885 ;
        RECT 677.795 1.195 678.125 1.525 ;
        RECT 677.795 -0.165 678.125 0.165 ;
        RECT 677.795 -1.525 678.125 -1.195 ;
        RECT 677.8 -1.525 678.12 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 679.155 7.995 679.485 8.325 ;
        RECT 679.155 2.555 679.485 2.885 ;
        RECT 679.155 1.195 679.485 1.525 ;
        RECT 679.155 -0.165 679.485 0.165 ;
        RECT 679.155 -1.525 679.485 -1.195 ;
        RECT 679.16 -1.525 679.48 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 680.515 7.995 680.845 8.325 ;
        RECT 680.515 2.555 680.845 2.885 ;
        RECT 680.515 1.195 680.845 1.525 ;
        RECT 680.515 -0.165 680.845 0.165 ;
        RECT 680.515 -1.525 680.845 -1.195 ;
        RECT 680.52 -1.525 680.84 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 681.875 7.995 682.205 8.325 ;
        RECT 681.875 2.555 682.205 2.885 ;
        RECT 681.875 1.195 682.205 1.525 ;
        RECT 681.875 -0.165 682.205 0.165 ;
        RECT 681.875 -1.525 682.205 -1.195 ;
        RECT 681.88 -1.525 682.2 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 683.235 7.995 683.565 8.325 ;
        RECT 683.235 2.555 683.565 2.885 ;
        RECT 683.235 1.195 683.565 1.525 ;
        RECT 683.235 -0.165 683.565 0.165 ;
        RECT 683.235 -1.525 683.565 -1.195 ;
        RECT 683.24 -1.525 683.56 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 684.595 7.995 684.925 8.325 ;
        RECT 684.595 2.555 684.925 2.885 ;
        RECT 684.595 1.195 684.925 1.525 ;
        RECT 684.595 -0.165 684.925 0.165 ;
        RECT 684.595 -1.525 684.925 -1.195 ;
        RECT 684.6 -1.525 684.92 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 685.955 7.995 686.285 8.325 ;
        RECT 685.955 2.555 686.285 2.885 ;
        RECT 685.955 1.195 686.285 1.525 ;
        RECT 685.955 -0.165 686.285 0.165 ;
        RECT 685.955 -1.525 686.285 -1.195 ;
        RECT 685.96 -1.525 686.28 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 687.315 7.995 687.645 8.325 ;
        RECT 687.315 2.555 687.645 2.885 ;
        RECT 687.315 1.195 687.645 1.525 ;
        RECT 687.315 -0.165 687.645 0.165 ;
        RECT 687.315 -1.525 687.645 -1.195 ;
        RECT 687.32 -1.525 687.64 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 688.675 7.995 689.005 8.325 ;
        RECT 688.675 2.555 689.005 2.885 ;
        RECT 688.675 1.195 689.005 1.525 ;
        RECT 688.675 -0.165 689.005 0.165 ;
        RECT 688.675 -1.525 689.005 -1.195 ;
        RECT 688.68 -1.525 689 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 690.035 7.995 690.365 8.325 ;
        RECT 690.035 2.555 690.365 2.885 ;
        RECT 690.035 1.195 690.365 1.525 ;
        RECT 690.035 -0.165 690.365 0.165 ;
        RECT 690.035 -1.525 690.365 -1.195 ;
        RECT 690.04 -1.525 690.36 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 691.395 7.995 691.725 8.325 ;
        RECT 691.395 2.555 691.725 2.885 ;
        RECT 691.395 1.195 691.725 1.525 ;
        RECT 691.395 -0.165 691.725 0.165 ;
        RECT 691.395 -1.525 691.725 -1.195 ;
        RECT 691.4 -1.525 691.72 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 692.755 7.995 693.085 8.325 ;
        RECT 692.755 2.555 693.085 2.885 ;
        RECT 692.755 1.195 693.085 1.525 ;
        RECT 692.755 -0.165 693.085 0.165 ;
        RECT 692.755 -1.525 693.085 -1.195 ;
        RECT 692.76 -1.525 693.08 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 694.115 7.995 694.445 8.325 ;
        RECT 694.115 2.555 694.445 2.885 ;
        RECT 694.115 1.195 694.445 1.525 ;
        RECT 694.115 -0.165 694.445 0.165 ;
        RECT 694.115 -1.525 694.445 -1.195 ;
        RECT 694.12 -1.525 694.44 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 695.475 7.995 695.805 8.325 ;
        RECT 695.475 2.555 695.805 2.885 ;
        RECT 695.475 1.195 695.805 1.525 ;
        RECT 695.475 -0.165 695.805 0.165 ;
        RECT 695.475 -1.525 695.805 -1.195 ;
        RECT 695.48 -1.525 695.8 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 696.835 7.995 697.165 8.325 ;
        RECT 696.835 2.555 697.165 2.885 ;
        RECT 696.835 1.195 697.165 1.525 ;
        RECT 696.835 -0.165 697.165 0.165 ;
        RECT 696.835 -1.525 697.165 -1.195 ;
        RECT 696.84 -1.525 697.16 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 698.195 7.995 698.525 8.325 ;
        RECT 698.195 2.555 698.525 2.885 ;
        RECT 698.195 1.195 698.525 1.525 ;
        RECT 698.195 -0.165 698.525 0.165 ;
        RECT 698.195 -1.525 698.525 -1.195 ;
        RECT 698.2 -1.525 698.52 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 699.555 7.995 699.885 8.325 ;
        RECT 699.555 2.555 699.885 2.885 ;
        RECT 699.555 1.195 699.885 1.525 ;
        RECT 699.555 -0.165 699.885 0.165 ;
        RECT 699.555 -1.525 699.885 -1.195 ;
        RECT 699.56 -1.525 699.88 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 700.915 7.995 701.245 8.325 ;
        RECT 700.915 2.555 701.245 2.885 ;
        RECT 700.915 1.195 701.245 1.525 ;
        RECT 700.915 -0.165 701.245 0.165 ;
        RECT 700.915 -1.525 701.245 -1.195 ;
        RECT 700.92 -1.525 701.24 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 702.275 7.995 702.605 8.325 ;
        RECT 702.275 2.555 702.605 2.885 ;
        RECT 702.275 1.195 702.605 1.525 ;
        RECT 702.275 -0.165 702.605 0.165 ;
        RECT 702.275 -1.525 702.605 -1.195 ;
        RECT 702.28 -1.525 702.6 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 703.635 7.995 703.965 8.325 ;
        RECT 703.635 2.555 703.965 2.885 ;
        RECT 703.635 1.195 703.965 1.525 ;
        RECT 703.635 -0.165 703.965 0.165 ;
        RECT 703.635 -1.525 703.965 -1.195 ;
        RECT 703.64 -1.525 703.96 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 704.995 7.995 705.325 8.325 ;
        RECT 704.995 2.555 705.325 2.885 ;
        RECT 704.995 1.195 705.325 1.525 ;
        RECT 704.995 -0.165 705.325 0.165 ;
        RECT 704.995 -1.525 705.325 -1.195 ;
        RECT 705 -1.525 705.32 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 706.355 7.995 706.685 8.325 ;
        RECT 706.355 2.555 706.685 2.885 ;
        RECT 706.355 1.195 706.685 1.525 ;
        RECT 706.355 -0.165 706.685 0.165 ;
        RECT 706.355 -1.525 706.685 -1.195 ;
        RECT 706.36 -1.525 706.68 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 707.715 7.995 708.045 8.325 ;
        RECT 707.715 2.555 708.045 2.885 ;
        RECT 707.715 1.195 708.045 1.525 ;
        RECT 707.715 -0.165 708.045 0.165 ;
        RECT 707.715 -1.525 708.045 -1.195 ;
        RECT 707.72 -1.525 708.04 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 709.075 7.995 709.405 8.325 ;
        RECT 709.075 2.555 709.405 2.885 ;
        RECT 709.075 1.195 709.405 1.525 ;
        RECT 709.075 -0.165 709.405 0.165 ;
        RECT 709.075 -1.525 709.405 -1.195 ;
        RECT 709.08 -1.525 709.4 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 710.435 7.995 710.765 8.325 ;
        RECT 710.435 2.555 710.765 2.885 ;
        RECT 710.435 1.195 710.765 1.525 ;
        RECT 710.435 -0.165 710.765 0.165 ;
        RECT 710.435 -1.525 710.765 -1.195 ;
        RECT 710.44 -1.525 710.76 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 711.795 7.995 712.125 8.325 ;
        RECT 711.795 2.555 712.125 2.885 ;
        RECT 711.795 1.195 712.125 1.525 ;
        RECT 711.795 -0.165 712.125 0.165 ;
        RECT 711.795 -1.525 712.125 -1.195 ;
        RECT 711.8 -1.525 712.12 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 713.155 7.995 713.485 8.325 ;
        RECT 713.155 2.555 713.485 2.885 ;
        RECT 713.155 1.195 713.485 1.525 ;
        RECT 713.155 -0.165 713.485 0.165 ;
        RECT 713.155 -1.525 713.485 -1.195 ;
        RECT 713.16 -1.525 713.48 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 714.515 7.995 714.845 8.325 ;
        RECT 714.515 2.555 714.845 2.885 ;
        RECT 714.515 1.195 714.845 1.525 ;
        RECT 714.515 -0.165 714.845 0.165 ;
        RECT 714.515 -1.525 714.845 -1.195 ;
        RECT 714.52 -1.525 714.84 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 715.875 7.995 716.205 8.325 ;
        RECT 715.875 2.555 716.205 2.885 ;
        RECT 715.875 1.195 716.205 1.525 ;
        RECT 715.875 -0.165 716.205 0.165 ;
        RECT 715.875 -1.525 716.205 -1.195 ;
        RECT 715.88 -1.525 716.2 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 717.235 7.995 717.565 8.325 ;
        RECT 717.235 2.555 717.565 2.885 ;
        RECT 717.235 1.195 717.565 1.525 ;
        RECT 717.235 -0.165 717.565 0.165 ;
        RECT 717.235 -1.525 717.565 -1.195 ;
        RECT 717.24 -1.525 717.56 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 718.595 7.995 718.925 8.325 ;
        RECT 718.595 2.555 718.925 2.885 ;
        RECT 718.595 1.195 718.925 1.525 ;
        RECT 718.595 -0.165 718.925 0.165 ;
        RECT 718.595 -1.525 718.925 -1.195 ;
        RECT 718.6 -1.525 718.92 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 719.955 7.995 720.285 8.325 ;
        RECT 719.955 2.555 720.285 2.885 ;
        RECT 719.955 1.195 720.285 1.525 ;
        RECT 719.955 -0.165 720.285 0.165 ;
        RECT 719.955 -1.525 720.285 -1.195 ;
        RECT 719.96 -1.525 720.28 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 721.315 7.995 721.645 8.325 ;
        RECT 721.315 2.555 721.645 2.885 ;
        RECT 721.315 1.195 721.645 1.525 ;
        RECT 721.315 -0.165 721.645 0.165 ;
        RECT 721.315 -1.525 721.645 -1.195 ;
        RECT 721.32 -1.525 721.64 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 722.675 7.995 723.005 8.325 ;
        RECT 722.675 2.555 723.005 2.885 ;
        RECT 722.675 1.195 723.005 1.525 ;
        RECT 722.675 -0.165 723.005 0.165 ;
        RECT 722.675 -1.525 723.005 -1.195 ;
        RECT 722.68 -1.525 723 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 724.035 7.995 724.365 8.325 ;
        RECT 724.035 2.555 724.365 2.885 ;
        RECT 724.035 1.195 724.365 1.525 ;
        RECT 724.035 -0.165 724.365 0.165 ;
        RECT 724.035 -1.525 724.365 -1.195 ;
        RECT 724.04 -1.525 724.36 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 725.395 7.995 725.725 8.325 ;
        RECT 725.395 2.555 725.725 2.885 ;
        RECT 725.395 1.195 725.725 1.525 ;
        RECT 725.395 -0.165 725.725 0.165 ;
        RECT 725.395 -1.525 725.725 -1.195 ;
        RECT 725.4 -1.525 725.72 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 726.755 7.995 727.085 8.325 ;
        RECT 726.755 2.555 727.085 2.885 ;
        RECT 726.755 1.195 727.085 1.525 ;
        RECT 726.755 -0.165 727.085 0.165 ;
        RECT 726.755 -1.525 727.085 -1.195 ;
        RECT 726.76 -1.525 727.08 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 728.115 7.995 728.445 8.325 ;
        RECT 728.115 2.555 728.445 2.885 ;
        RECT 728.115 1.195 728.445 1.525 ;
        RECT 728.115 -0.165 728.445 0.165 ;
        RECT 728.115 -1.525 728.445 -1.195 ;
        RECT 728.12 -1.525 728.44 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 729.475 7.995 729.805 8.325 ;
        RECT 729.475 2.555 729.805 2.885 ;
        RECT 729.475 1.195 729.805 1.525 ;
        RECT 729.475 -0.165 729.805 0.165 ;
        RECT 729.475 -1.525 729.805 -1.195 ;
        RECT 729.48 -1.525 729.8 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 730.835 7.995 731.165 8.325 ;
        RECT 730.835 2.555 731.165 2.885 ;
        RECT 730.835 1.195 731.165 1.525 ;
        RECT 730.835 -0.165 731.165 0.165 ;
        RECT 730.835 -1.525 731.165 -1.195 ;
        RECT 730.84 -1.525 731.16 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 732.195 7.995 732.525 8.325 ;
        RECT 732.195 2.555 732.525 2.885 ;
        RECT 732.195 1.195 732.525 1.525 ;
        RECT 732.195 -0.165 732.525 0.165 ;
        RECT 732.195 -1.525 732.525 -1.195 ;
        RECT 732.2 -1.525 732.52 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 733.555 7.995 733.885 8.325 ;
        RECT 733.555 2.555 733.885 2.885 ;
        RECT 733.555 1.195 733.885 1.525 ;
        RECT 733.555 -0.165 733.885 0.165 ;
        RECT 733.555 -1.525 733.885 -1.195 ;
        RECT 733.56 -1.525 733.88 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 734.915 7.995 735.245 8.325 ;
        RECT 734.915 2.555 735.245 2.885 ;
        RECT 734.915 1.195 735.245 1.525 ;
        RECT 734.915 -0.165 735.245 0.165 ;
        RECT 734.915 -1.525 735.245 -1.195 ;
        RECT 734.92 -1.525 735.24 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 736.275 7.995 736.605 8.325 ;
        RECT 736.275 2.555 736.605 2.885 ;
        RECT 736.275 1.195 736.605 1.525 ;
        RECT 736.275 -0.165 736.605 0.165 ;
        RECT 736.275 -1.525 736.605 -1.195 ;
        RECT 736.28 -1.525 736.6 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 737.635 7.995 737.965 8.325 ;
        RECT 737.635 2.555 737.965 2.885 ;
        RECT 737.635 1.195 737.965 1.525 ;
        RECT 737.635 -0.165 737.965 0.165 ;
        RECT 737.635 -1.525 737.965 -1.195 ;
        RECT 737.64 -1.525 737.96 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 738.995 7.995 739.325 8.325 ;
        RECT 738.995 2.555 739.325 2.885 ;
        RECT 738.995 1.195 739.325 1.525 ;
        RECT 738.995 -0.165 739.325 0.165 ;
        RECT 738.995 -1.525 739.325 -1.195 ;
        RECT 739 -1.525 739.32 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 740.355 7.995 740.685 8.325 ;
        RECT 740.355 2.555 740.685 2.885 ;
        RECT 740.355 1.195 740.685 1.525 ;
        RECT 740.355 -0.165 740.685 0.165 ;
        RECT 740.355 -1.525 740.685 -1.195 ;
        RECT 740.36 -1.525 740.68 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 741.715 7.995 742.045 8.325 ;
        RECT 741.715 2.555 742.045 2.885 ;
        RECT 741.715 1.195 742.045 1.525 ;
        RECT 741.715 -0.165 742.045 0.165 ;
        RECT 741.715 -1.525 742.045 -1.195 ;
        RECT 741.72 -1.525 742.04 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 743.075 7.995 743.405 8.325 ;
        RECT 743.075 2.555 743.405 2.885 ;
        RECT 743.075 1.195 743.405 1.525 ;
        RECT 743.075 -0.165 743.405 0.165 ;
        RECT 743.075 -1.525 743.405 -1.195 ;
        RECT 743.08 -1.525 743.4 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 744.435 7.995 744.765 8.325 ;
        RECT 744.435 2.555 744.765 2.885 ;
        RECT 744.435 1.195 744.765 1.525 ;
        RECT 744.435 -0.165 744.765 0.165 ;
        RECT 744.435 -1.525 744.765 -1.195 ;
        RECT 744.44 -1.525 744.76 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 745.795 7.995 746.125 8.325 ;
        RECT 745.795 2.555 746.125 2.885 ;
        RECT 745.795 1.195 746.125 1.525 ;
        RECT 745.795 -0.165 746.125 0.165 ;
        RECT 745.795 -1.525 746.125 -1.195 ;
        RECT 745.8 -1.525 746.12 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 747.155 7.995 747.485 8.325 ;
        RECT 747.155 2.555 747.485 2.885 ;
        RECT 747.155 1.195 747.485 1.525 ;
        RECT 747.155 -0.165 747.485 0.165 ;
        RECT 747.155 -1.525 747.485 -1.195 ;
        RECT 747.16 -1.525 747.48 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 748.515 7.995 748.845 8.325 ;
        RECT 748.515 2.555 748.845 2.885 ;
        RECT 748.515 1.195 748.845 1.525 ;
        RECT 748.515 -0.165 748.845 0.165 ;
        RECT 748.515 -1.525 748.845 -1.195 ;
        RECT 748.52 -1.525 748.84 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 749.875 7.995 750.205 8.325 ;
        RECT 749.875 2.555 750.205 2.885 ;
        RECT 749.875 1.195 750.205 1.525 ;
        RECT 749.875 -0.165 750.205 0.165 ;
        RECT 749.875 -1.525 750.205 -1.195 ;
        RECT 749.88 -1.525 750.2 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 751.235 7.995 751.565 8.325 ;
        RECT 751.235 2.555 751.565 2.885 ;
        RECT 751.235 1.195 751.565 1.525 ;
        RECT 751.235 -0.165 751.565 0.165 ;
        RECT 751.235 -1.525 751.565 -1.195 ;
        RECT 751.24 -1.525 751.56 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 752.595 7.995 752.925 8.325 ;
        RECT 752.595 2.555 752.925 2.885 ;
        RECT 752.595 1.195 752.925 1.525 ;
        RECT 752.595 -0.165 752.925 0.165 ;
        RECT 752.595 -1.525 752.925 -1.195 ;
        RECT 752.6 -1.525 752.92 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 753.955 7.995 754.285 8.325 ;
        RECT 753.955 2.555 754.285 2.885 ;
        RECT 753.955 1.195 754.285 1.525 ;
        RECT 753.955 -0.165 754.285 0.165 ;
        RECT 753.955 -1.525 754.285 -1.195 ;
        RECT 753.96 -1.525 754.28 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 755.315 7.995 755.645 8.325 ;
        RECT 755.315 2.555 755.645 2.885 ;
        RECT 755.315 1.195 755.645 1.525 ;
        RECT 755.315 -0.165 755.645 0.165 ;
        RECT 755.315 -1.525 755.645 -1.195 ;
        RECT 755.32 -1.525 755.64 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 756.675 7.995 757.005 8.325 ;
        RECT 756.675 2.555 757.005 2.885 ;
        RECT 756.675 1.195 757.005 1.525 ;
        RECT 756.675 -0.165 757.005 0.165 ;
        RECT 756.675 -1.525 757.005 -1.195 ;
        RECT 756.68 -1.525 757 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 758.035 7.995 758.365 8.325 ;
        RECT 758.035 2.555 758.365 2.885 ;
        RECT 758.035 1.195 758.365 1.525 ;
        RECT 758.035 -0.165 758.365 0.165 ;
        RECT 758.035 -1.525 758.365 -1.195 ;
        RECT 758.04 -1.525 758.36 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 759.395 7.995 759.725 8.325 ;
        RECT 759.395 2.555 759.725 2.885 ;
        RECT 759.395 1.195 759.725 1.525 ;
        RECT 759.395 -0.165 759.725 0.165 ;
        RECT 759.395 -1.525 759.725 -1.195 ;
        RECT 759.4 -1.525 759.72 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 760.755 7.995 761.085 8.325 ;
        RECT 760.755 2.555 761.085 2.885 ;
        RECT 760.755 1.195 761.085 1.525 ;
        RECT 760.755 -0.165 761.085 0.165 ;
        RECT 760.755 -1.525 761.085 -1.195 ;
        RECT 760.76 -1.525 761.08 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 762.115 7.995 762.445 8.325 ;
        RECT 762.115 2.555 762.445 2.885 ;
        RECT 762.115 1.195 762.445 1.525 ;
        RECT 762.115 -0.165 762.445 0.165 ;
        RECT 762.115 -1.525 762.445 -1.195 ;
        RECT 762.12 -1.525 762.44 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 763.475 7.995 763.805 8.325 ;
        RECT 763.475 5.275 763.805 5.605 ;
        RECT 763.475 2.555 763.805 2.885 ;
        RECT 763.475 1.195 763.805 1.525 ;
        RECT 763.475 -0.165 763.805 0.165 ;
        RECT 763.475 -1.525 763.805 -1.195 ;
        RECT 763.48 -1.525 763.8 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 764.835 7.995 765.165 8.325 ;
        RECT 764.835 5.275 765.165 5.605 ;
        RECT 764.835 3.915 765.165 4.245 ;
        RECT 764.835 2.555 765.165 2.885 ;
        RECT 764.835 1.195 765.165 1.525 ;
        RECT 764.835 -0.165 765.165 0.165 ;
        RECT 764.835 -1.525 765.165 -1.195 ;
        RECT 764.84 -1.525 765.16 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 766.195 7.995 766.525 8.325 ;
        RECT 766.195 5.275 766.525 5.605 ;
        RECT 766.195 3.915 766.525 4.245 ;
        RECT 766.195 2.555 766.525 2.885 ;
        RECT 766.195 1.195 766.525 1.525 ;
        RECT 766.195 -0.165 766.525 0.165 ;
        RECT 766.195 -1.525 766.525 -1.195 ;
        RECT 766.2 -1.525 766.52 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 767.555 7.995 767.885 8.325 ;
        RECT 767.555 6.635 767.885 6.965 ;
        RECT 767.555 5.275 767.885 5.605 ;
        RECT 767.555 3.915 767.885 4.245 ;
        RECT 767.555 2.555 767.885 2.885 ;
        RECT 767.555 1.195 767.885 1.525 ;
        RECT 767.555 -0.165 767.885 0.165 ;
        RECT 767.555 -1.525 767.885 -1.195 ;
        RECT 767.56 -1.525 767.88 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 768.915 7.995 769.245 8.325 ;
        RECT 768.915 6.635 769.245 6.965 ;
        RECT 768.915 5.275 769.245 5.605 ;
        RECT 768.915 3.915 769.245 4.245 ;
        RECT 768.915 2.555 769.245 2.885 ;
        RECT 768.915 1.195 769.245 1.525 ;
        RECT 768.915 -0.165 769.245 0.165 ;
        RECT 768.915 -1.525 769.245 -1.195 ;
        RECT 768.92 -1.525 769.24 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 320.115 7.995 320.445 8.325 ;
        RECT 320.115 2.555 320.445 2.885 ;
        RECT 320.115 1.195 320.445 1.525 ;
        RECT 320.115 -0.165 320.445 0.165 ;
        RECT 320.115 -1.525 320.445 -1.195 ;
        RECT 320.12 -1.525 320.44 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 321.475 7.995 321.805 8.325 ;
        RECT 321.475 2.555 321.805 2.885 ;
        RECT 321.475 1.195 321.805 1.525 ;
        RECT 321.475 -0.165 321.805 0.165 ;
        RECT 321.475 -1.525 321.805 -1.195 ;
        RECT 321.48 -1.525 321.8 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 322.835 7.995 323.165 8.325 ;
        RECT 322.835 2.555 323.165 2.885 ;
        RECT 322.835 1.195 323.165 1.525 ;
        RECT 322.835 -0.165 323.165 0.165 ;
        RECT 322.835 -1.525 323.165 -1.195 ;
        RECT 322.84 -1.525 323.16 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.195 7.995 324.525 8.325 ;
        RECT 324.195 2.555 324.525 2.885 ;
        RECT 324.195 1.195 324.525 1.525 ;
        RECT 324.195 -0.165 324.525 0.165 ;
        RECT 324.195 -1.525 324.525 -1.195 ;
        RECT 324.2 -1.525 324.52 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 325.555 7.995 325.885 8.325 ;
        RECT 325.555 2.555 325.885 2.885 ;
        RECT 325.555 1.195 325.885 1.525 ;
        RECT 325.555 -0.165 325.885 0.165 ;
        RECT 325.555 -1.525 325.885 -1.195 ;
        RECT 325.56 -1.525 325.88 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 326.915 7.995 327.245 8.325 ;
        RECT 326.915 2.555 327.245 2.885 ;
        RECT 326.915 1.195 327.245 1.525 ;
        RECT 326.915 -0.165 327.245 0.165 ;
        RECT 326.915 -1.525 327.245 -1.195 ;
        RECT 326.92 -1.525 327.24 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 328.275 7.995 328.605 8.325 ;
        RECT 328.275 2.555 328.605 2.885 ;
        RECT 328.275 1.195 328.605 1.525 ;
        RECT 328.275 -0.165 328.605 0.165 ;
        RECT 328.275 -1.525 328.605 -1.195 ;
        RECT 328.28 -1.525 328.6 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 329.635 7.995 329.965 8.325 ;
        RECT 329.635 2.555 329.965 2.885 ;
        RECT 329.635 1.195 329.965 1.525 ;
        RECT 329.635 -0.165 329.965 0.165 ;
        RECT 329.635 -1.525 329.965 -1.195 ;
        RECT 329.64 -1.525 329.96 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.995 7.995 331.325 8.325 ;
        RECT 330.995 2.555 331.325 2.885 ;
        RECT 330.995 1.195 331.325 1.525 ;
        RECT 330.995 -0.165 331.325 0.165 ;
        RECT 330.995 -1.525 331.325 -1.195 ;
        RECT 331 -1.525 331.32 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 332.355 7.995 332.685 8.325 ;
        RECT 332.355 2.555 332.685 2.885 ;
        RECT 332.355 1.195 332.685 1.525 ;
        RECT 332.355 -0.165 332.685 0.165 ;
        RECT 332.355 -1.525 332.685 -1.195 ;
        RECT 332.36 -1.525 332.68 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 333.715 7.995 334.045 8.325 ;
        RECT 333.715 2.555 334.045 2.885 ;
        RECT 333.715 1.195 334.045 1.525 ;
        RECT 333.715 -0.165 334.045 0.165 ;
        RECT 333.715 -1.525 334.045 -1.195 ;
        RECT 333.72 -1.525 334.04 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.075 7.995 335.405 8.325 ;
        RECT 335.075 2.555 335.405 2.885 ;
        RECT 335.075 1.195 335.405 1.525 ;
        RECT 335.075 -0.165 335.405 0.165 ;
        RECT 335.075 -1.525 335.405 -1.195 ;
        RECT 335.08 -1.525 335.4 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 336.435 7.995 336.765 8.325 ;
        RECT 336.435 2.555 336.765 2.885 ;
        RECT 336.435 1.195 336.765 1.525 ;
        RECT 336.435 -0.165 336.765 0.165 ;
        RECT 336.435 -1.525 336.765 -1.195 ;
        RECT 336.44 -1.525 336.76 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 337.795 7.995 338.125 8.325 ;
        RECT 337.795 2.555 338.125 2.885 ;
        RECT 337.795 1.195 338.125 1.525 ;
        RECT 337.795 -0.165 338.125 0.165 ;
        RECT 337.795 -1.525 338.125 -1.195 ;
        RECT 337.8 -1.525 338.12 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 339.155 7.995 339.485 8.325 ;
        RECT 339.155 2.555 339.485 2.885 ;
        RECT 339.155 1.195 339.485 1.525 ;
        RECT 339.155 -0.165 339.485 0.165 ;
        RECT 339.155 -1.525 339.485 -1.195 ;
        RECT 339.16 -1.525 339.48 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 340.515 7.995 340.845 8.325 ;
        RECT 340.515 2.555 340.845 2.885 ;
        RECT 340.515 1.195 340.845 1.525 ;
        RECT 340.515 -0.165 340.845 0.165 ;
        RECT 340.515 -1.525 340.845 -1.195 ;
        RECT 340.52 -1.525 340.84 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 341.875 7.995 342.205 8.325 ;
        RECT 341.875 2.555 342.205 2.885 ;
        RECT 341.875 1.195 342.205 1.525 ;
        RECT 341.875 -0.165 342.205 0.165 ;
        RECT 341.875 -1.525 342.205 -1.195 ;
        RECT 341.88 -1.525 342.2 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 343.235 7.995 343.565 8.325 ;
        RECT 343.235 2.555 343.565 2.885 ;
        RECT 343.235 1.195 343.565 1.525 ;
        RECT 343.235 -0.165 343.565 0.165 ;
        RECT 343.235 -1.525 343.565 -1.195 ;
        RECT 343.24 -1.525 343.56 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 344.595 7.995 344.925 8.325 ;
        RECT 344.595 2.555 344.925 2.885 ;
        RECT 344.595 1.195 344.925 1.525 ;
        RECT 344.595 -0.165 344.925 0.165 ;
        RECT 344.595 -1.525 344.925 -1.195 ;
        RECT 344.6 -1.525 344.92 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 345.955 7.995 346.285 8.325 ;
        RECT 345.955 2.555 346.285 2.885 ;
        RECT 345.955 1.195 346.285 1.525 ;
        RECT 345.955 -0.165 346.285 0.165 ;
        RECT 345.955 -1.525 346.285 -1.195 ;
        RECT 345.96 -1.525 346.28 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 347.315 7.995 347.645 8.325 ;
        RECT 347.315 2.555 347.645 2.885 ;
        RECT 347.315 1.195 347.645 1.525 ;
        RECT 347.315 -0.165 347.645 0.165 ;
        RECT 347.315 -1.525 347.645 -1.195 ;
        RECT 347.32 -1.525 347.64 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 348.675 7.995 349.005 8.325 ;
        RECT 348.675 2.555 349.005 2.885 ;
        RECT 348.675 1.195 349.005 1.525 ;
        RECT 348.675 -0.165 349.005 0.165 ;
        RECT 348.675 -1.525 349.005 -1.195 ;
        RECT 348.68 -1.525 349 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 350.035 7.995 350.365 8.325 ;
        RECT 350.035 2.555 350.365 2.885 ;
        RECT 350.035 1.195 350.365 1.525 ;
        RECT 350.035 -0.165 350.365 0.165 ;
        RECT 350.035 -1.525 350.365 -1.195 ;
        RECT 350.04 -1.525 350.36 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 351.395 7.995 351.725 8.325 ;
        RECT 351.395 2.555 351.725 2.885 ;
        RECT 351.395 1.195 351.725 1.525 ;
        RECT 351.395 -0.165 351.725 0.165 ;
        RECT 351.395 -1.525 351.725 -1.195 ;
        RECT 351.4 -1.525 351.72 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 352.755 7.995 353.085 8.325 ;
        RECT 352.755 2.555 353.085 2.885 ;
        RECT 352.755 1.195 353.085 1.525 ;
        RECT 352.755 -0.165 353.085 0.165 ;
        RECT 352.755 -1.525 353.085 -1.195 ;
        RECT 352.76 -1.525 353.08 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.115 7.995 354.445 8.325 ;
        RECT 354.115 2.555 354.445 2.885 ;
        RECT 354.115 1.195 354.445 1.525 ;
        RECT 354.115 -0.165 354.445 0.165 ;
        RECT 354.115 -1.525 354.445 -1.195 ;
        RECT 354.12 -1.525 354.44 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 355.475 7.995 355.805 8.325 ;
        RECT 355.475 2.555 355.805 2.885 ;
        RECT 355.475 1.195 355.805 1.525 ;
        RECT 355.475 -0.165 355.805 0.165 ;
        RECT 355.475 -1.525 355.805 -1.195 ;
        RECT 355.48 -1.525 355.8 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 356.835 7.995 357.165 8.325 ;
        RECT 356.835 2.555 357.165 2.885 ;
        RECT 356.835 1.195 357.165 1.525 ;
        RECT 356.835 -0.165 357.165 0.165 ;
        RECT 356.835 -1.525 357.165 -1.195 ;
        RECT 356.84 -1.525 357.16 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 358.195 7.995 358.525 8.325 ;
        RECT 358.195 2.555 358.525 2.885 ;
        RECT 358.195 1.195 358.525 1.525 ;
        RECT 358.195 -0.165 358.525 0.165 ;
        RECT 358.195 -1.525 358.525 -1.195 ;
        RECT 358.2 -1.525 358.52 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 359.555 7.995 359.885 8.325 ;
        RECT 359.555 2.555 359.885 2.885 ;
        RECT 359.555 1.195 359.885 1.525 ;
        RECT 359.555 -0.165 359.885 0.165 ;
        RECT 359.555 -1.525 359.885 -1.195 ;
        RECT 359.56 -1.525 359.88 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 360.915 7.995 361.245 8.325 ;
        RECT 360.915 2.555 361.245 2.885 ;
        RECT 360.915 1.195 361.245 1.525 ;
        RECT 360.915 -0.165 361.245 0.165 ;
        RECT 360.915 -1.525 361.245 -1.195 ;
        RECT 360.92 -1.525 361.24 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 362.275 7.995 362.605 8.325 ;
        RECT 362.275 2.555 362.605 2.885 ;
        RECT 362.275 1.195 362.605 1.525 ;
        RECT 362.275 -0.165 362.605 0.165 ;
        RECT 362.275 -1.525 362.605 -1.195 ;
        RECT 362.28 -1.525 362.6 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 363.635 7.995 363.965 8.325 ;
        RECT 363.635 2.555 363.965 2.885 ;
        RECT 363.635 1.195 363.965 1.525 ;
        RECT 363.635 -0.165 363.965 0.165 ;
        RECT 363.635 -1.525 363.965 -1.195 ;
        RECT 363.64 -1.525 363.96 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 364.995 7.995 365.325 8.325 ;
        RECT 364.995 2.555 365.325 2.885 ;
        RECT 364.995 1.195 365.325 1.525 ;
        RECT 364.995 -0.165 365.325 0.165 ;
        RECT 364.995 -1.525 365.325 -1.195 ;
        RECT 365 -1.525 365.32 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 366.355 7.995 366.685 8.325 ;
        RECT 366.355 2.555 366.685 2.885 ;
        RECT 366.355 1.195 366.685 1.525 ;
        RECT 366.355 -0.165 366.685 0.165 ;
        RECT 366.355 -1.525 366.685 -1.195 ;
        RECT 366.36 -1.525 366.68 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 367.715 7.995 368.045 8.325 ;
        RECT 367.715 2.555 368.045 2.885 ;
        RECT 367.715 1.195 368.045 1.525 ;
        RECT 367.715 -0.165 368.045 0.165 ;
        RECT 367.715 -1.525 368.045 -1.195 ;
        RECT 367.72 -1.525 368.04 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 369.075 7.995 369.405 8.325 ;
        RECT 369.075 2.555 369.405 2.885 ;
        RECT 369.075 1.195 369.405 1.525 ;
        RECT 369.075 -0.165 369.405 0.165 ;
        RECT 369.075 -1.525 369.405 -1.195 ;
        RECT 369.08 -1.525 369.4 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 370.435 7.995 370.765 8.325 ;
        RECT 370.435 2.555 370.765 2.885 ;
        RECT 370.435 1.195 370.765 1.525 ;
        RECT 370.435 -0.165 370.765 0.165 ;
        RECT 370.435 -1.525 370.765 -1.195 ;
        RECT 370.44 -1.525 370.76 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 371.795 7.995 372.125 8.325 ;
        RECT 371.795 2.555 372.125 2.885 ;
        RECT 371.795 1.195 372.125 1.525 ;
        RECT 371.795 -0.165 372.125 0.165 ;
        RECT 371.795 -1.525 372.125 -1.195 ;
        RECT 371.8 -1.525 372.12 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 373.155 7.995 373.485 8.325 ;
        RECT 373.155 2.555 373.485 2.885 ;
        RECT 373.155 1.195 373.485 1.525 ;
        RECT 373.155 -0.165 373.485 0.165 ;
        RECT 373.155 -1.525 373.485 -1.195 ;
        RECT 373.16 -1.525 373.48 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 374.515 7.995 374.845 8.325 ;
        RECT 374.515 2.555 374.845 2.885 ;
        RECT 374.515 1.195 374.845 1.525 ;
        RECT 374.515 -0.165 374.845 0.165 ;
        RECT 374.515 -1.525 374.845 -1.195 ;
        RECT 374.52 -1.525 374.84 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 375.875 7.995 376.205 8.325 ;
        RECT 375.875 2.555 376.205 2.885 ;
        RECT 375.875 1.195 376.205 1.525 ;
        RECT 375.875 -0.165 376.205 0.165 ;
        RECT 375.875 -1.525 376.205 -1.195 ;
        RECT 375.88 -1.525 376.2 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 377.235 7.995 377.565 8.325 ;
        RECT 377.235 2.555 377.565 2.885 ;
        RECT 377.235 1.195 377.565 1.525 ;
        RECT 377.235 -0.165 377.565 0.165 ;
        RECT 377.235 -1.525 377.565 -1.195 ;
        RECT 377.24 -1.525 377.56 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 378.595 7.995 378.925 8.325 ;
        RECT 378.595 2.555 378.925 2.885 ;
        RECT 378.595 1.195 378.925 1.525 ;
        RECT 378.595 -0.165 378.925 0.165 ;
        RECT 378.595 -1.525 378.925 -1.195 ;
        RECT 378.6 -1.525 378.92 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 379.955 7.995 380.285 8.325 ;
        RECT 379.955 2.555 380.285 2.885 ;
        RECT 379.955 1.195 380.285 1.525 ;
        RECT 379.955 -0.165 380.285 0.165 ;
        RECT 379.955 -1.525 380.285 -1.195 ;
        RECT 379.96 -1.525 380.28 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 381.315 7.995 381.645 8.325 ;
        RECT 381.315 2.555 381.645 2.885 ;
        RECT 381.315 1.195 381.645 1.525 ;
        RECT 381.315 -0.165 381.645 0.165 ;
        RECT 381.315 -1.525 381.645 -1.195 ;
        RECT 381.32 -1.525 381.64 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 382.675 7.995 383.005 8.325 ;
        RECT 382.675 2.555 383.005 2.885 ;
        RECT 382.675 1.195 383.005 1.525 ;
        RECT 382.675 -0.165 383.005 0.165 ;
        RECT 382.675 -1.525 383.005 -1.195 ;
        RECT 382.68 -1.525 383 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 384.035 7.995 384.365 8.325 ;
        RECT 384.035 2.555 384.365 2.885 ;
        RECT 384.035 1.195 384.365 1.525 ;
        RECT 384.035 -0.165 384.365 0.165 ;
        RECT 384.035 -1.525 384.365 -1.195 ;
        RECT 384.04 -1.525 384.36 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 385.395 7.995 385.725 8.325 ;
        RECT 385.395 2.555 385.725 2.885 ;
        RECT 385.395 1.195 385.725 1.525 ;
        RECT 385.395 -0.165 385.725 0.165 ;
        RECT 385.395 -1.525 385.725 -1.195 ;
        RECT 385.4 -1.525 385.72 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 386.755 7.995 387.085 8.325 ;
        RECT 386.755 2.555 387.085 2.885 ;
        RECT 386.755 1.195 387.085 1.525 ;
        RECT 386.755 -0.165 387.085 0.165 ;
        RECT 386.755 -1.525 387.085 -1.195 ;
        RECT 386.76 -1.525 387.08 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 388.115 7.995 388.445 8.325 ;
        RECT 388.115 2.555 388.445 2.885 ;
        RECT 388.115 1.195 388.445 1.525 ;
        RECT 388.115 -0.165 388.445 0.165 ;
        RECT 388.115 -1.525 388.445 -1.195 ;
        RECT 388.12 -1.525 388.44 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 389.475 7.995 389.805 8.325 ;
        RECT 389.475 2.555 389.805 2.885 ;
        RECT 389.475 1.195 389.805 1.525 ;
        RECT 389.475 -0.165 389.805 0.165 ;
        RECT 389.475 -1.525 389.805 -1.195 ;
        RECT 389.48 -1.525 389.8 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 390.835 7.995 391.165 8.325 ;
        RECT 390.835 2.555 391.165 2.885 ;
        RECT 390.835 1.195 391.165 1.525 ;
        RECT 390.835 -0.165 391.165 0.165 ;
        RECT 390.835 -1.525 391.165 -1.195 ;
        RECT 390.84 -1.525 391.16 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 392.195 7.995 392.525 8.325 ;
        RECT 392.195 2.555 392.525 2.885 ;
        RECT 392.195 1.195 392.525 1.525 ;
        RECT 392.195 -0.165 392.525 0.165 ;
        RECT 392.195 -1.525 392.525 -1.195 ;
        RECT 392.2 -1.525 392.52 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 393.555 7.995 393.885 8.325 ;
        RECT 393.555 2.555 393.885 2.885 ;
        RECT 393.555 1.195 393.885 1.525 ;
        RECT 393.555 -0.165 393.885 0.165 ;
        RECT 393.555 -1.525 393.885 -1.195 ;
        RECT 393.56 -1.525 393.88 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 394.915 7.995 395.245 8.325 ;
        RECT 394.915 2.555 395.245 2.885 ;
        RECT 394.915 1.195 395.245 1.525 ;
        RECT 394.915 -0.165 395.245 0.165 ;
        RECT 394.915 -1.525 395.245 -1.195 ;
        RECT 394.92 -1.525 395.24 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 396.275 7.995 396.605 8.325 ;
        RECT 396.275 2.555 396.605 2.885 ;
        RECT 396.275 1.195 396.605 1.525 ;
        RECT 396.275 -0.165 396.605 0.165 ;
        RECT 396.275 -1.525 396.605 -1.195 ;
        RECT 396.28 -1.525 396.6 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 397.635 7.995 397.965 8.325 ;
        RECT 397.635 2.555 397.965 2.885 ;
        RECT 397.635 1.195 397.965 1.525 ;
        RECT 397.635 -0.165 397.965 0.165 ;
        RECT 397.635 -1.525 397.965 -1.195 ;
        RECT 397.64 -1.525 397.96 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 398.995 7.995 399.325 8.325 ;
        RECT 398.995 2.555 399.325 2.885 ;
        RECT 398.995 1.195 399.325 1.525 ;
        RECT 398.995 -0.165 399.325 0.165 ;
        RECT 398.995 -1.525 399.325 -1.195 ;
        RECT 399 -1.525 399.32 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 400.355 7.995 400.685 8.325 ;
        RECT 400.355 2.555 400.685 2.885 ;
        RECT 400.355 1.195 400.685 1.525 ;
        RECT 400.355 -0.165 400.685 0.165 ;
        RECT 400.355 -1.525 400.685 -1.195 ;
        RECT 400.36 -1.525 400.68 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 401.715 7.995 402.045 8.325 ;
        RECT 401.715 2.555 402.045 2.885 ;
        RECT 401.715 1.195 402.045 1.525 ;
        RECT 401.715 -0.165 402.045 0.165 ;
        RECT 401.715 -1.525 402.045 -1.195 ;
        RECT 401.72 -1.525 402.04 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 403.075 7.995 403.405 8.325 ;
        RECT 403.075 2.555 403.405 2.885 ;
        RECT 403.075 1.195 403.405 1.525 ;
        RECT 403.075 -0.165 403.405 0.165 ;
        RECT 403.075 -1.525 403.405 -1.195 ;
        RECT 403.08 -1.525 403.4 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 404.435 7.995 404.765 8.325 ;
        RECT 404.435 2.555 404.765 2.885 ;
        RECT 404.435 1.195 404.765 1.525 ;
        RECT 404.435 -0.165 404.765 0.165 ;
        RECT 404.435 -1.525 404.765 -1.195 ;
        RECT 404.44 -1.525 404.76 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 405.795 7.995 406.125 8.325 ;
        RECT 405.795 2.555 406.125 2.885 ;
        RECT 405.795 1.195 406.125 1.525 ;
        RECT 405.795 -0.165 406.125 0.165 ;
        RECT 405.795 -1.525 406.125 -1.195 ;
        RECT 405.8 -1.525 406.12 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 407.155 7.995 407.485 8.325 ;
        RECT 407.155 2.555 407.485 2.885 ;
        RECT 407.155 1.195 407.485 1.525 ;
        RECT 407.155 -0.165 407.485 0.165 ;
        RECT 407.155 -1.525 407.485 -1.195 ;
        RECT 407.16 -1.525 407.48 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 408.515 7.995 408.845 8.325 ;
        RECT 408.515 2.555 408.845 2.885 ;
        RECT 408.515 1.195 408.845 1.525 ;
        RECT 408.515 -0.165 408.845 0.165 ;
        RECT 408.515 -1.525 408.845 -1.195 ;
        RECT 408.52 -1.525 408.84 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 409.875 7.995 410.205 8.325 ;
        RECT 409.875 2.555 410.205 2.885 ;
        RECT 409.875 1.195 410.205 1.525 ;
        RECT 409.875 -0.165 410.205 0.165 ;
        RECT 409.875 -1.525 410.205 -1.195 ;
        RECT 409.88 -1.525 410.2 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 411.235 7.995 411.565 8.325 ;
        RECT 411.235 2.555 411.565 2.885 ;
        RECT 411.235 1.195 411.565 1.525 ;
        RECT 411.235 -0.165 411.565 0.165 ;
        RECT 411.235 -1.525 411.565 -1.195 ;
        RECT 411.24 -1.525 411.56 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 412.595 7.995 412.925 8.325 ;
        RECT 412.595 2.555 412.925 2.885 ;
        RECT 412.595 1.195 412.925 1.525 ;
        RECT 412.595 -0.165 412.925 0.165 ;
        RECT 412.595 -1.525 412.925 -1.195 ;
        RECT 412.6 -1.525 412.92 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 413.955 7.995 414.285 8.325 ;
        RECT 413.955 2.555 414.285 2.885 ;
        RECT 413.955 1.195 414.285 1.525 ;
        RECT 413.955 -0.165 414.285 0.165 ;
        RECT 413.955 -1.525 414.285 -1.195 ;
        RECT 413.96 -1.525 414.28 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 415.315 7.995 415.645 8.325 ;
        RECT 415.315 2.555 415.645 2.885 ;
        RECT 415.315 1.195 415.645 1.525 ;
        RECT 415.315 -0.165 415.645 0.165 ;
        RECT 415.315 -1.525 415.645 -1.195 ;
        RECT 415.32 -1.525 415.64 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 416.675 7.995 417.005 8.325 ;
        RECT 416.675 2.555 417.005 2.885 ;
        RECT 416.675 1.195 417.005 1.525 ;
        RECT 416.675 -0.165 417.005 0.165 ;
        RECT 416.675 -1.525 417.005 -1.195 ;
        RECT 416.68 -1.525 417 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 418.035 7.995 418.365 8.325 ;
        RECT 418.035 2.555 418.365 2.885 ;
        RECT 418.035 1.195 418.365 1.525 ;
        RECT 418.035 -0.165 418.365 0.165 ;
        RECT 418.035 -1.525 418.365 -1.195 ;
        RECT 418.04 -1.525 418.36 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 419.395 7.995 419.725 8.325 ;
        RECT 419.395 2.555 419.725 2.885 ;
        RECT 419.395 1.195 419.725 1.525 ;
        RECT 419.395 -0.165 419.725 0.165 ;
        RECT 419.395 -1.525 419.725 -1.195 ;
        RECT 419.4 -1.525 419.72 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 420.755 7.995 421.085 8.325 ;
        RECT 420.755 2.555 421.085 2.885 ;
        RECT 420.755 1.195 421.085 1.525 ;
        RECT 420.755 -0.165 421.085 0.165 ;
        RECT 420.755 -1.525 421.085 -1.195 ;
        RECT 420.76 -1.525 421.08 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 422.115 7.995 422.445 8.325 ;
        RECT 422.115 2.555 422.445 2.885 ;
        RECT 422.115 1.195 422.445 1.525 ;
        RECT 422.115 -0.165 422.445 0.165 ;
        RECT 422.115 -1.525 422.445 -1.195 ;
        RECT 422.12 -1.525 422.44 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 423.475 7.995 423.805 8.325 ;
        RECT 423.475 2.555 423.805 2.885 ;
        RECT 423.475 1.195 423.805 1.525 ;
        RECT 423.475 -0.165 423.805 0.165 ;
        RECT 423.475 -1.525 423.805 -1.195 ;
        RECT 423.48 -1.525 423.8 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 424.835 7.995 425.165 8.325 ;
        RECT 424.835 2.555 425.165 2.885 ;
        RECT 424.835 1.195 425.165 1.525 ;
        RECT 424.835 -0.165 425.165 0.165 ;
        RECT 424.835 -1.525 425.165 -1.195 ;
        RECT 424.84 -1.525 425.16 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 426.195 7.995 426.525 8.325 ;
        RECT 426.195 2.555 426.525 2.885 ;
        RECT 426.195 1.195 426.525 1.525 ;
        RECT 426.195 -0.165 426.525 0.165 ;
        RECT 426.195 -1.525 426.525 -1.195 ;
        RECT 426.2 -1.525 426.52 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 427.555 7.995 427.885 8.325 ;
        RECT 427.555 2.555 427.885 2.885 ;
        RECT 427.555 1.195 427.885 1.525 ;
        RECT 427.555 -0.165 427.885 0.165 ;
        RECT 427.555 -1.525 427.885 -1.195 ;
        RECT 427.56 -1.525 427.88 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 428.915 7.995 429.245 8.325 ;
        RECT 428.915 2.555 429.245 2.885 ;
        RECT 428.915 1.195 429.245 1.525 ;
        RECT 428.915 -0.165 429.245 0.165 ;
        RECT 428.915 -1.525 429.245 -1.195 ;
        RECT 428.92 -1.525 429.24 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 430.275 7.995 430.605 8.325 ;
        RECT 430.275 2.555 430.605 2.885 ;
        RECT 430.275 1.195 430.605 1.525 ;
        RECT 430.275 -0.165 430.605 0.165 ;
        RECT 430.275 -1.525 430.605 -1.195 ;
        RECT 430.28 -1.525 430.6 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 431.635 7.995 431.965 8.325 ;
        RECT 431.635 2.555 431.965 2.885 ;
        RECT 431.635 1.195 431.965 1.525 ;
        RECT 431.635 -0.165 431.965 0.165 ;
        RECT 431.635 -1.525 431.965 -1.195 ;
        RECT 431.64 -1.525 431.96 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 432.995 7.995 433.325 8.325 ;
        RECT 432.995 2.555 433.325 2.885 ;
        RECT 432.995 1.195 433.325 1.525 ;
        RECT 432.995 -0.165 433.325 0.165 ;
        RECT 432.995 -1.525 433.325 -1.195 ;
        RECT 433 -1.525 433.32 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 434.355 7.995 434.685 8.325 ;
        RECT 434.355 2.555 434.685 2.885 ;
        RECT 434.355 1.195 434.685 1.525 ;
        RECT 434.355 -0.165 434.685 0.165 ;
        RECT 434.355 -1.525 434.685 -1.195 ;
        RECT 434.36 -1.525 434.68 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 435.715 7.995 436.045 8.325 ;
        RECT 435.715 2.555 436.045 2.885 ;
        RECT 435.715 1.195 436.045 1.525 ;
        RECT 435.715 -0.165 436.045 0.165 ;
        RECT 435.715 -1.525 436.045 -1.195 ;
        RECT 435.72 -1.525 436.04 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 437.075 7.995 437.405 8.325 ;
        RECT 437.075 2.555 437.405 2.885 ;
        RECT 437.075 1.195 437.405 1.525 ;
        RECT 437.075 -0.165 437.405 0.165 ;
        RECT 437.075 -1.525 437.405 -1.195 ;
        RECT 437.08 -1.525 437.4 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 438.435 7.995 438.765 8.325 ;
        RECT 438.435 2.555 438.765 2.885 ;
        RECT 438.435 1.195 438.765 1.525 ;
        RECT 438.435 -0.165 438.765 0.165 ;
        RECT 438.435 -1.525 438.765 -1.195 ;
        RECT 438.44 -1.525 438.76 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 439.795 7.995 440.125 8.325 ;
        RECT 439.795 2.555 440.125 2.885 ;
        RECT 439.795 1.195 440.125 1.525 ;
        RECT 439.795 -0.165 440.125 0.165 ;
        RECT 439.795 -1.525 440.125 -1.195 ;
        RECT 439.8 -1.525 440.12 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 441.155 7.995 441.485 8.325 ;
        RECT 441.155 2.555 441.485 2.885 ;
        RECT 441.155 1.195 441.485 1.525 ;
        RECT 441.155 -0.165 441.485 0.165 ;
        RECT 441.155 -1.525 441.485 -1.195 ;
        RECT 441.16 -1.525 441.48 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 442.515 7.995 442.845 8.325 ;
        RECT 442.515 2.555 442.845 2.885 ;
        RECT 442.515 1.195 442.845 1.525 ;
        RECT 442.515 -0.165 442.845 0.165 ;
        RECT 442.515 -1.525 442.845 -1.195 ;
        RECT 442.52 -1.525 442.84 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 443.875 7.995 444.205 8.325 ;
        RECT 443.875 2.555 444.205 2.885 ;
        RECT 443.875 1.195 444.205 1.525 ;
        RECT 443.875 -0.165 444.205 0.165 ;
        RECT 443.875 -1.525 444.205 -1.195 ;
        RECT 443.88 -1.525 444.2 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 445.235 7.995 445.565 8.325 ;
        RECT 445.235 2.555 445.565 2.885 ;
        RECT 445.235 1.195 445.565 1.525 ;
        RECT 445.235 -0.165 445.565 0.165 ;
        RECT 445.235 -1.525 445.565 -1.195 ;
        RECT 445.24 -1.525 445.56 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 446.595 7.995 446.925 8.325 ;
        RECT 446.595 2.555 446.925 2.885 ;
        RECT 446.595 1.195 446.925 1.525 ;
        RECT 446.595 -0.165 446.925 0.165 ;
        RECT 446.595 -1.525 446.925 -1.195 ;
        RECT 446.6 -1.525 446.92 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 447.955 7.995 448.285 8.325 ;
        RECT 447.955 2.555 448.285 2.885 ;
        RECT 447.955 1.195 448.285 1.525 ;
        RECT 447.955 -0.165 448.285 0.165 ;
        RECT 447.955 -1.525 448.285 -1.195 ;
        RECT 447.96 -1.525 448.28 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 449.315 7.995 449.645 8.325 ;
        RECT 449.315 2.555 449.645 2.885 ;
        RECT 449.315 1.195 449.645 1.525 ;
        RECT 449.315 -0.165 449.645 0.165 ;
        RECT 449.315 -1.525 449.645 -1.195 ;
        RECT 449.32 -1.525 449.64 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 450.675 7.995 451.005 8.325 ;
        RECT 450.675 2.555 451.005 2.885 ;
        RECT 450.675 1.195 451.005 1.525 ;
        RECT 450.675 -0.165 451.005 0.165 ;
        RECT 450.675 -1.525 451.005 -1.195 ;
        RECT 450.68 -1.525 451 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 452.035 7.995 452.365 8.325 ;
        RECT 452.035 2.555 452.365 2.885 ;
        RECT 452.035 1.195 452.365 1.525 ;
        RECT 452.035 -0.165 452.365 0.165 ;
        RECT 452.035 -1.525 452.365 -1.195 ;
        RECT 452.04 -1.525 452.36 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 453.395 7.995 453.725 8.325 ;
        RECT 453.395 2.555 453.725 2.885 ;
        RECT 453.395 1.195 453.725 1.525 ;
        RECT 453.395 -0.165 453.725 0.165 ;
        RECT 453.395 -1.525 453.725 -1.195 ;
        RECT 453.4 -1.525 453.72 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 454.755 7.995 455.085 8.325 ;
        RECT 454.755 2.555 455.085 2.885 ;
        RECT 454.755 1.195 455.085 1.525 ;
        RECT 454.755 -0.165 455.085 0.165 ;
        RECT 454.755 -1.525 455.085 -1.195 ;
        RECT 454.76 -1.525 455.08 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 456.115 7.995 456.445 8.325 ;
        RECT 456.115 2.555 456.445 2.885 ;
        RECT 456.115 1.195 456.445 1.525 ;
        RECT 456.115 -0.165 456.445 0.165 ;
        RECT 456.115 -1.525 456.445 -1.195 ;
        RECT 456.12 -1.525 456.44 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 457.475 7.995 457.805 8.325 ;
        RECT 457.475 2.555 457.805 2.885 ;
        RECT 457.475 1.195 457.805 1.525 ;
        RECT 457.475 -0.165 457.805 0.165 ;
        RECT 457.475 -1.525 457.805 -1.195 ;
        RECT 457.48 -1.525 457.8 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 458.835 7.995 459.165 8.325 ;
        RECT 458.835 2.555 459.165 2.885 ;
        RECT 458.835 1.195 459.165 1.525 ;
        RECT 458.835 -0.165 459.165 0.165 ;
        RECT 458.835 -1.525 459.165 -1.195 ;
        RECT 458.84 -1.525 459.16 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 460.195 7.995 460.525 8.325 ;
        RECT 460.195 2.555 460.525 2.885 ;
        RECT 460.195 1.195 460.525 1.525 ;
        RECT 460.195 -0.165 460.525 0.165 ;
        RECT 460.195 -1.525 460.525 -1.195 ;
        RECT 460.2 -1.525 460.52 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 461.555 7.995 461.885 8.325 ;
        RECT 461.555 2.555 461.885 2.885 ;
        RECT 461.555 1.195 461.885 1.525 ;
        RECT 461.555 -0.165 461.885 0.165 ;
        RECT 461.555 -1.525 461.885 -1.195 ;
        RECT 461.56 -1.525 461.88 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 462.915 7.995 463.245 8.325 ;
        RECT 462.915 2.555 463.245 2.885 ;
        RECT 462.915 1.195 463.245 1.525 ;
        RECT 462.915 -0.165 463.245 0.165 ;
        RECT 462.915 -1.525 463.245 -1.195 ;
        RECT 462.92 -1.525 463.24 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 464.275 7.995 464.605 8.325 ;
        RECT 464.275 2.555 464.605 2.885 ;
        RECT 464.275 1.195 464.605 1.525 ;
        RECT 464.275 -0.165 464.605 0.165 ;
        RECT 464.275 -1.525 464.605 -1.195 ;
        RECT 464.28 -1.525 464.6 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 465.635 7.995 465.965 8.325 ;
        RECT 465.635 2.555 465.965 2.885 ;
        RECT 465.635 1.195 465.965 1.525 ;
        RECT 465.635 -0.165 465.965 0.165 ;
        RECT 465.635 -1.525 465.965 -1.195 ;
        RECT 465.64 -1.525 465.96 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 466.995 7.995 467.325 8.325 ;
        RECT 466.995 2.555 467.325 2.885 ;
        RECT 466.995 1.195 467.325 1.525 ;
        RECT 466.995 -0.165 467.325 0.165 ;
        RECT 466.995 -1.525 467.325 -1.195 ;
        RECT 467 -1.525 467.32 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 468.355 7.995 468.685 8.325 ;
        RECT 468.355 2.555 468.685 2.885 ;
        RECT 468.355 1.195 468.685 1.525 ;
        RECT 468.355 -0.165 468.685 0.165 ;
        RECT 468.355 -1.525 468.685 -1.195 ;
        RECT 468.36 -1.525 468.68 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 469.715 7.995 470.045 8.325 ;
        RECT 469.715 2.555 470.045 2.885 ;
        RECT 469.715 1.195 470.045 1.525 ;
        RECT 469.715 -0.165 470.045 0.165 ;
        RECT 469.715 -1.525 470.045 -1.195 ;
        RECT 469.72 -1.525 470.04 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 471.075 7.995 471.405 8.325 ;
        RECT 471.075 2.555 471.405 2.885 ;
        RECT 471.075 1.195 471.405 1.525 ;
        RECT 471.075 -0.165 471.405 0.165 ;
        RECT 471.075 -1.525 471.405 -1.195 ;
        RECT 471.08 -1.525 471.4 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 472.435 7.995 472.765 8.325 ;
        RECT 472.435 2.555 472.765 2.885 ;
        RECT 472.435 1.195 472.765 1.525 ;
        RECT 472.435 -0.165 472.765 0.165 ;
        RECT 472.435 -1.525 472.765 -1.195 ;
        RECT 472.44 -1.525 472.76 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 473.795 7.995 474.125 8.325 ;
        RECT 473.795 2.555 474.125 2.885 ;
        RECT 473.795 1.195 474.125 1.525 ;
        RECT 473.795 -0.165 474.125 0.165 ;
        RECT 473.795 -1.525 474.125 -1.195 ;
        RECT 473.8 -1.525 474.12 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 475.155 7.995 475.485 8.325 ;
        RECT 475.155 2.555 475.485 2.885 ;
        RECT 475.155 1.195 475.485 1.525 ;
        RECT 475.155 -0.165 475.485 0.165 ;
        RECT 475.155 -1.525 475.485 -1.195 ;
        RECT 475.16 -1.525 475.48 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 476.515 7.995 476.845 8.325 ;
        RECT 476.515 2.555 476.845 2.885 ;
        RECT 476.515 1.195 476.845 1.525 ;
        RECT 476.515 -0.165 476.845 0.165 ;
        RECT 476.515 -1.525 476.845 -1.195 ;
        RECT 476.52 -1.525 476.84 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 477.875 7.995 478.205 8.325 ;
        RECT 477.875 2.555 478.205 2.885 ;
        RECT 477.875 1.195 478.205 1.525 ;
        RECT 477.875 -0.165 478.205 0.165 ;
        RECT 477.875 -1.525 478.205 -1.195 ;
        RECT 477.88 -1.525 478.2 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 479.235 7.995 479.565 8.325 ;
        RECT 479.235 2.555 479.565 2.885 ;
        RECT 479.235 1.195 479.565 1.525 ;
        RECT 479.235 -0.165 479.565 0.165 ;
        RECT 479.235 -1.525 479.565 -1.195 ;
        RECT 479.24 -1.525 479.56 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 480.595 7.995 480.925 8.325 ;
        RECT 480.595 2.555 480.925 2.885 ;
        RECT 480.595 1.195 480.925 1.525 ;
        RECT 480.595 -0.165 480.925 0.165 ;
        RECT 480.595 -1.525 480.925 -1.195 ;
        RECT 480.6 -1.525 480.92 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 481.955 7.995 482.285 8.325 ;
        RECT 481.955 2.555 482.285 2.885 ;
        RECT 481.955 1.195 482.285 1.525 ;
        RECT 481.955 -0.165 482.285 0.165 ;
        RECT 481.955 -1.525 482.285 -1.195 ;
        RECT 481.96 -1.525 482.28 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 483.315 7.995 483.645 8.325 ;
        RECT 483.315 2.555 483.645 2.885 ;
        RECT 483.315 1.195 483.645 1.525 ;
        RECT 483.315 -0.165 483.645 0.165 ;
        RECT 483.315 -1.525 483.645 -1.195 ;
        RECT 483.32 -1.525 483.64 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 484.675 7.995 485.005 8.325 ;
        RECT 484.675 2.555 485.005 2.885 ;
        RECT 484.675 1.195 485.005 1.525 ;
        RECT 484.675 -0.165 485.005 0.165 ;
        RECT 484.675 -1.525 485.005 -1.195 ;
        RECT 484.68 -1.525 485 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 486.035 7.995 486.365 8.325 ;
        RECT 486.035 2.555 486.365 2.885 ;
        RECT 486.035 1.195 486.365 1.525 ;
        RECT 486.035 -0.165 486.365 0.165 ;
        RECT 486.035 -1.525 486.365 -1.195 ;
        RECT 486.04 -1.525 486.36 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 487.395 7.995 487.725 8.325 ;
        RECT 487.395 2.555 487.725 2.885 ;
        RECT 487.395 1.195 487.725 1.525 ;
        RECT 487.395 -0.165 487.725 0.165 ;
        RECT 487.395 -1.525 487.725 -1.195 ;
        RECT 487.4 -1.525 487.72 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 488.755 7.995 489.085 8.325 ;
        RECT 488.755 2.555 489.085 2.885 ;
        RECT 488.755 1.195 489.085 1.525 ;
        RECT 488.755 -0.165 489.085 0.165 ;
        RECT 488.755 -1.525 489.085 -1.195 ;
        RECT 488.76 -1.525 489.08 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 490.115 7.995 490.445 8.325 ;
        RECT 490.115 2.555 490.445 2.885 ;
        RECT 490.115 1.195 490.445 1.525 ;
        RECT 490.115 -0.165 490.445 0.165 ;
        RECT 490.115 -1.525 490.445 -1.195 ;
        RECT 490.12 -1.525 490.44 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 491.475 7.995 491.805 8.325 ;
        RECT 491.475 2.555 491.805 2.885 ;
        RECT 491.475 1.195 491.805 1.525 ;
        RECT 491.475 -0.165 491.805 0.165 ;
        RECT 491.475 -1.525 491.805 -1.195 ;
        RECT 491.48 -1.525 491.8 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 492.835 7.995 493.165 8.325 ;
        RECT 492.835 2.555 493.165 2.885 ;
        RECT 492.835 1.195 493.165 1.525 ;
        RECT 492.835 -0.165 493.165 0.165 ;
        RECT 492.835 -1.525 493.165 -1.195 ;
        RECT 492.84 -1.525 493.16 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 494.195 7.995 494.525 8.325 ;
        RECT 494.195 2.555 494.525 2.885 ;
        RECT 494.195 1.195 494.525 1.525 ;
        RECT 494.195 -0.165 494.525 0.165 ;
        RECT 494.195 -1.525 494.525 -1.195 ;
        RECT 494.2 -1.525 494.52 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 495.555 7.995 495.885 8.325 ;
        RECT 495.555 2.555 495.885 2.885 ;
        RECT 495.555 1.195 495.885 1.525 ;
        RECT 495.555 -0.165 495.885 0.165 ;
        RECT 495.555 -1.525 495.885 -1.195 ;
        RECT 495.56 -1.525 495.88 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 496.915 7.995 497.245 8.325 ;
        RECT 496.915 2.555 497.245 2.885 ;
        RECT 496.915 1.195 497.245 1.525 ;
        RECT 496.915 -0.165 497.245 0.165 ;
        RECT 496.915 -1.525 497.245 -1.195 ;
        RECT 496.92 -1.525 497.24 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 498.275 7.995 498.605 8.325 ;
        RECT 498.275 2.555 498.605 2.885 ;
        RECT 498.275 1.195 498.605 1.525 ;
        RECT 498.275 -0.165 498.605 0.165 ;
        RECT 498.275 -1.525 498.605 -1.195 ;
        RECT 498.28 -1.525 498.6 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 499.635 7.995 499.965 8.325 ;
        RECT 499.635 2.555 499.965 2.885 ;
        RECT 499.635 1.195 499.965 1.525 ;
        RECT 499.635 -0.165 499.965 0.165 ;
        RECT 499.635 -1.525 499.965 -1.195 ;
        RECT 499.64 -1.525 499.96 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 500.995 7.995 501.325 8.325 ;
        RECT 500.995 2.555 501.325 2.885 ;
        RECT 500.995 1.195 501.325 1.525 ;
        RECT 500.995 -0.165 501.325 0.165 ;
        RECT 500.995 -1.525 501.325 -1.195 ;
        RECT 501 -1.525 501.32 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 502.355 7.995 502.685 8.325 ;
        RECT 502.355 2.555 502.685 2.885 ;
        RECT 502.355 1.195 502.685 1.525 ;
        RECT 502.355 -0.165 502.685 0.165 ;
        RECT 502.355 -1.525 502.685 -1.195 ;
        RECT 502.36 -1.525 502.68 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 503.715 7.995 504.045 8.325 ;
        RECT 503.715 2.555 504.045 2.885 ;
        RECT 503.715 1.195 504.045 1.525 ;
        RECT 503.715 -0.165 504.045 0.165 ;
        RECT 503.715 -1.525 504.045 -1.195 ;
        RECT 503.72 -1.525 504.04 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 505.075 7.995 505.405 8.325 ;
        RECT 505.075 2.555 505.405 2.885 ;
        RECT 505.075 1.195 505.405 1.525 ;
        RECT 505.075 -0.165 505.405 0.165 ;
        RECT 505.075 -1.525 505.405 -1.195 ;
        RECT 505.08 -1.525 505.4 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 506.435 7.995 506.765 8.325 ;
        RECT 506.435 2.555 506.765 2.885 ;
        RECT 506.435 1.195 506.765 1.525 ;
        RECT 506.435 -0.165 506.765 0.165 ;
        RECT 506.435 -1.525 506.765 -1.195 ;
        RECT 506.44 -1.525 506.76 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 507.795 7.995 508.125 8.325 ;
        RECT 507.795 2.555 508.125 2.885 ;
        RECT 507.795 1.195 508.125 1.525 ;
        RECT 507.795 -0.165 508.125 0.165 ;
        RECT 507.795 -1.525 508.125 -1.195 ;
        RECT 507.8 -1.525 508.12 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 509.155 7.995 509.485 8.325 ;
        RECT 509.155 2.555 509.485 2.885 ;
        RECT 509.155 1.195 509.485 1.525 ;
        RECT 509.155 -0.165 509.485 0.165 ;
        RECT 509.155 -1.525 509.485 -1.195 ;
        RECT 509.16 -1.525 509.48 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 510.515 7.995 510.845 8.325 ;
        RECT 510.515 2.555 510.845 2.885 ;
        RECT 510.515 1.195 510.845 1.525 ;
        RECT 510.515 -0.165 510.845 0.165 ;
        RECT 510.515 -1.525 510.845 -1.195 ;
        RECT 510.52 -1.525 510.84 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 511.875 7.995 512.205 8.325 ;
        RECT 511.875 2.555 512.205 2.885 ;
        RECT 511.875 1.195 512.205 1.525 ;
        RECT 511.875 -0.165 512.205 0.165 ;
        RECT 511.875 -1.525 512.205 -1.195 ;
        RECT 511.88 -1.525 512.2 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 513.235 7.995 513.565 8.325 ;
        RECT 513.235 2.555 513.565 2.885 ;
        RECT 513.235 1.195 513.565 1.525 ;
        RECT 513.235 -0.165 513.565 0.165 ;
        RECT 513.235 -1.525 513.565 -1.195 ;
        RECT 513.24 -1.525 513.56 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 514.595 7.995 514.925 8.325 ;
        RECT 514.595 2.555 514.925 2.885 ;
        RECT 514.595 1.195 514.925 1.525 ;
        RECT 514.595 -0.165 514.925 0.165 ;
        RECT 514.595 -1.525 514.925 -1.195 ;
        RECT 514.6 -1.525 514.92 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 515.955 7.995 516.285 8.325 ;
        RECT 515.955 2.555 516.285 2.885 ;
        RECT 515.955 1.195 516.285 1.525 ;
        RECT 515.955 -0.165 516.285 0.165 ;
        RECT 515.955 -1.525 516.285 -1.195 ;
        RECT 515.96 -1.525 516.28 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 517.315 7.995 517.645 8.325 ;
        RECT 517.315 2.555 517.645 2.885 ;
        RECT 517.315 1.195 517.645 1.525 ;
        RECT 517.315 -0.165 517.645 0.165 ;
        RECT 517.315 -1.525 517.645 -1.195 ;
        RECT 517.32 -1.525 517.64 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 518.675 7.995 519.005 8.325 ;
        RECT 518.675 2.555 519.005 2.885 ;
        RECT 518.675 1.195 519.005 1.525 ;
        RECT 518.675 -0.165 519.005 0.165 ;
        RECT 518.675 -1.525 519.005 -1.195 ;
        RECT 518.68 -1.525 519 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 520.035 7.995 520.365 8.325 ;
        RECT 520.035 2.555 520.365 2.885 ;
        RECT 520.035 1.195 520.365 1.525 ;
        RECT 520.035 -0.165 520.365 0.165 ;
        RECT 520.035 -1.525 520.365 -1.195 ;
        RECT 520.04 -1.525 520.36 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 521.395 7.995 521.725 8.325 ;
        RECT 521.395 2.555 521.725 2.885 ;
        RECT 521.395 1.195 521.725 1.525 ;
        RECT 521.395 -0.165 521.725 0.165 ;
        RECT 521.395 -1.525 521.725 -1.195 ;
        RECT 521.4 -1.525 521.72 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 522.755 7.995 523.085 8.325 ;
        RECT 522.755 2.555 523.085 2.885 ;
        RECT 522.755 1.195 523.085 1.525 ;
        RECT 522.755 -0.165 523.085 0.165 ;
        RECT 522.755 -1.525 523.085 -1.195 ;
        RECT 522.76 -1.525 523.08 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 524.115 7.995 524.445 8.325 ;
        RECT 524.115 2.555 524.445 2.885 ;
        RECT 524.115 1.195 524.445 1.525 ;
        RECT 524.115 -0.165 524.445 0.165 ;
        RECT 524.115 -1.525 524.445 -1.195 ;
        RECT 524.12 -1.525 524.44 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 525.475 7.995 525.805 8.325 ;
        RECT 525.475 2.555 525.805 2.885 ;
        RECT 525.475 1.195 525.805 1.525 ;
        RECT 525.475 -0.165 525.805 0.165 ;
        RECT 525.475 -1.525 525.805 -1.195 ;
        RECT 525.48 -1.525 525.8 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 526.835 7.995 527.165 8.325 ;
        RECT 526.835 2.555 527.165 2.885 ;
        RECT 526.835 1.195 527.165 1.525 ;
        RECT 526.835 -0.165 527.165 0.165 ;
        RECT 526.835 -1.525 527.165 -1.195 ;
        RECT 526.84 -1.525 527.16 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 528.195 7.995 528.525 8.325 ;
        RECT 528.195 2.555 528.525 2.885 ;
        RECT 528.195 1.195 528.525 1.525 ;
        RECT 528.195 -0.165 528.525 0.165 ;
        RECT 528.195 -1.525 528.525 -1.195 ;
        RECT 528.2 -1.525 528.52 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 529.555 7.995 529.885 8.325 ;
        RECT 529.555 2.555 529.885 2.885 ;
        RECT 529.555 1.195 529.885 1.525 ;
        RECT 529.555 -0.165 529.885 0.165 ;
        RECT 529.555 -1.525 529.885 -1.195 ;
        RECT 529.56 -1.525 529.88 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 530.915 7.995 531.245 8.325 ;
        RECT 530.915 2.555 531.245 2.885 ;
        RECT 530.915 1.195 531.245 1.525 ;
        RECT 530.915 -0.165 531.245 0.165 ;
        RECT 530.915 -1.525 531.245 -1.195 ;
        RECT 530.92 -1.525 531.24 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 532.275 7.995 532.605 8.325 ;
        RECT 532.275 2.555 532.605 2.885 ;
        RECT 532.275 1.195 532.605 1.525 ;
        RECT 532.275 -0.165 532.605 0.165 ;
        RECT 532.275 -1.525 532.605 -1.195 ;
        RECT 532.28 -1.525 532.6 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 533.635 7.995 533.965 8.325 ;
        RECT 533.635 2.555 533.965 2.885 ;
        RECT 533.635 1.195 533.965 1.525 ;
        RECT 533.635 -0.165 533.965 0.165 ;
        RECT 533.635 -1.525 533.965 -1.195 ;
        RECT 533.64 -1.525 533.96 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 534.995 7.995 535.325 8.325 ;
        RECT 534.995 2.555 535.325 2.885 ;
        RECT 534.995 1.195 535.325 1.525 ;
        RECT 534.995 -0.165 535.325 0.165 ;
        RECT 534.995 -1.525 535.325 -1.195 ;
        RECT 535 -1.525 535.32 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 536.355 7.995 536.685 8.325 ;
        RECT 536.355 2.555 536.685 2.885 ;
        RECT 536.355 1.195 536.685 1.525 ;
        RECT 536.355 -0.165 536.685 0.165 ;
        RECT 536.355 -1.525 536.685 -1.195 ;
        RECT 536.36 -1.525 536.68 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 537.715 7.995 538.045 8.325 ;
        RECT 537.715 2.555 538.045 2.885 ;
        RECT 537.715 1.195 538.045 1.525 ;
        RECT 537.715 -0.165 538.045 0.165 ;
        RECT 537.715 -1.525 538.045 -1.195 ;
        RECT 537.72 -1.525 538.04 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 539.075 7.995 539.405 8.325 ;
        RECT 539.075 2.555 539.405 2.885 ;
        RECT 539.075 1.195 539.405 1.525 ;
        RECT 539.075 -0.165 539.405 0.165 ;
        RECT 539.075 -1.525 539.405 -1.195 ;
        RECT 539.08 -1.525 539.4 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 540.435 7.995 540.765 8.325 ;
        RECT 540.435 2.555 540.765 2.885 ;
        RECT 540.435 1.195 540.765 1.525 ;
        RECT 540.435 -0.165 540.765 0.165 ;
        RECT 540.435 -1.525 540.765 -1.195 ;
        RECT 540.44 -1.525 540.76 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 541.795 7.995 542.125 8.325 ;
        RECT 541.795 2.555 542.125 2.885 ;
        RECT 541.795 1.195 542.125 1.525 ;
        RECT 541.795 -0.165 542.125 0.165 ;
        RECT 541.795 -1.525 542.125 -1.195 ;
        RECT 541.8 -1.525 542.12 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 543.155 7.995 543.485 8.325 ;
        RECT 543.155 2.555 543.485 2.885 ;
        RECT 543.155 1.195 543.485 1.525 ;
        RECT 543.155 -0.165 543.485 0.165 ;
        RECT 543.155 -1.525 543.485 -1.195 ;
        RECT 543.16 -1.525 543.48 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 544.515 7.995 544.845 8.325 ;
        RECT 544.515 2.555 544.845 2.885 ;
        RECT 544.515 1.195 544.845 1.525 ;
        RECT 544.515 -0.165 544.845 0.165 ;
        RECT 544.515 -1.525 544.845 -1.195 ;
        RECT 544.52 -1.525 544.84 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 545.88 -1.525 546.2 9 ;
        RECT 545.875 7.995 546.205 8.325 ;
        RECT 545.875 2.555 546.205 2.885 ;
        RECT 545.875 1.195 546.205 1.525 ;
        RECT 545.875 -0.165 546.205 0.165 ;
        RECT 545.875 -1.525 546.205 -1.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.995 7.995 93.325 8.325 ;
        RECT 92.995 2.555 93.325 2.885 ;
        RECT 92.995 1.195 93.325 1.525 ;
        RECT 92.995 -0.165 93.325 0.165 ;
        RECT 92.995 -1.525 93.325 -1.195 ;
        RECT 93 -1.525 93.32 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.355 7.995 94.685 8.325 ;
        RECT 94.355 2.555 94.685 2.885 ;
        RECT 94.355 1.195 94.685 1.525 ;
        RECT 94.355 -0.165 94.685 0.165 ;
        RECT 94.355 -1.525 94.685 -1.195 ;
        RECT 94.36 -1.525 94.68 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.715 7.995 96.045 8.325 ;
        RECT 95.715 2.555 96.045 2.885 ;
        RECT 95.715 1.195 96.045 1.525 ;
        RECT 95.715 -0.165 96.045 0.165 ;
        RECT 95.715 -1.525 96.045 -1.195 ;
        RECT 95.72 -1.525 96.04 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.075 7.995 97.405 8.325 ;
        RECT 97.075 2.555 97.405 2.885 ;
        RECT 97.075 1.195 97.405 1.525 ;
        RECT 97.075 -0.165 97.405 0.165 ;
        RECT 97.075 -1.525 97.405 -1.195 ;
        RECT 97.08 -1.525 97.4 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.435 7.995 98.765 8.325 ;
        RECT 98.435 2.555 98.765 2.885 ;
        RECT 98.435 1.195 98.765 1.525 ;
        RECT 98.435 -0.165 98.765 0.165 ;
        RECT 98.435 -1.525 98.765 -1.195 ;
        RECT 98.44 -1.525 98.76 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.795 7.995 100.125 8.325 ;
        RECT 99.795 2.555 100.125 2.885 ;
        RECT 99.795 1.195 100.125 1.525 ;
        RECT 99.795 -0.165 100.125 0.165 ;
        RECT 99.795 -1.525 100.125 -1.195 ;
        RECT 99.8 -1.525 100.12 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.155 7.995 101.485 8.325 ;
        RECT 101.155 2.555 101.485 2.885 ;
        RECT 101.155 1.195 101.485 1.525 ;
        RECT 101.155 -0.165 101.485 0.165 ;
        RECT 101.155 -1.525 101.485 -1.195 ;
        RECT 101.16 -1.525 101.48 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.515 7.995 102.845 8.325 ;
        RECT 102.515 2.555 102.845 2.885 ;
        RECT 102.515 1.195 102.845 1.525 ;
        RECT 102.515 -0.165 102.845 0.165 ;
        RECT 102.515 -1.525 102.845 -1.195 ;
        RECT 102.52 -1.525 102.84 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.875 7.995 104.205 8.325 ;
        RECT 103.875 2.555 104.205 2.885 ;
        RECT 103.875 1.195 104.205 1.525 ;
        RECT 103.875 -0.165 104.205 0.165 ;
        RECT 103.875 -1.525 104.205 -1.195 ;
        RECT 103.88 -1.525 104.2 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.235 7.995 105.565 8.325 ;
        RECT 105.235 2.555 105.565 2.885 ;
        RECT 105.235 1.195 105.565 1.525 ;
        RECT 105.235 -0.165 105.565 0.165 ;
        RECT 105.235 -1.525 105.565 -1.195 ;
        RECT 105.24 -1.525 105.56 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.595 7.995 106.925 8.325 ;
        RECT 106.595 2.555 106.925 2.885 ;
        RECT 106.595 1.195 106.925 1.525 ;
        RECT 106.595 -0.165 106.925 0.165 ;
        RECT 106.595 -1.525 106.925 -1.195 ;
        RECT 106.6 -1.525 106.92 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.955 7.995 108.285 8.325 ;
        RECT 107.955 2.555 108.285 2.885 ;
        RECT 107.955 1.195 108.285 1.525 ;
        RECT 107.955 -0.165 108.285 0.165 ;
        RECT 107.955 -1.525 108.285 -1.195 ;
        RECT 107.96 -1.525 108.28 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.315 7.995 109.645 8.325 ;
        RECT 109.315 2.555 109.645 2.885 ;
        RECT 109.315 1.195 109.645 1.525 ;
        RECT 109.315 -0.165 109.645 0.165 ;
        RECT 109.315 -1.525 109.645 -1.195 ;
        RECT 109.32 -1.525 109.64 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.675 7.995 111.005 8.325 ;
        RECT 110.675 2.555 111.005 2.885 ;
        RECT 110.675 1.195 111.005 1.525 ;
        RECT 110.675 -0.165 111.005 0.165 ;
        RECT 110.675 -1.525 111.005 -1.195 ;
        RECT 110.68 -1.525 111 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.035 7.995 112.365 8.325 ;
        RECT 112.035 2.555 112.365 2.885 ;
        RECT 112.035 1.195 112.365 1.525 ;
        RECT 112.035 -0.165 112.365 0.165 ;
        RECT 112.035 -1.525 112.365 -1.195 ;
        RECT 112.04 -1.525 112.36 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.395 7.995 113.725 8.325 ;
        RECT 113.395 2.555 113.725 2.885 ;
        RECT 113.395 1.195 113.725 1.525 ;
        RECT 113.395 -0.165 113.725 0.165 ;
        RECT 113.395 -1.525 113.725 -1.195 ;
        RECT 113.4 -1.525 113.72 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.755 7.995 115.085 8.325 ;
        RECT 114.755 2.555 115.085 2.885 ;
        RECT 114.755 1.195 115.085 1.525 ;
        RECT 114.755 -0.165 115.085 0.165 ;
        RECT 114.755 -1.525 115.085 -1.195 ;
        RECT 114.76 -1.525 115.08 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.115 7.995 116.445 8.325 ;
        RECT 116.115 2.555 116.445 2.885 ;
        RECT 116.115 1.195 116.445 1.525 ;
        RECT 116.115 -0.165 116.445 0.165 ;
        RECT 116.115 -1.525 116.445 -1.195 ;
        RECT 116.12 -1.525 116.44 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 117.475 7.995 117.805 8.325 ;
        RECT 117.475 2.555 117.805 2.885 ;
        RECT 117.475 1.195 117.805 1.525 ;
        RECT 117.475 -0.165 117.805 0.165 ;
        RECT 117.475 -1.525 117.805 -1.195 ;
        RECT 117.48 -1.525 117.8 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.835 7.995 119.165 8.325 ;
        RECT 118.835 2.555 119.165 2.885 ;
        RECT 118.835 1.195 119.165 1.525 ;
        RECT 118.835 -0.165 119.165 0.165 ;
        RECT 118.835 -1.525 119.165 -1.195 ;
        RECT 118.84 -1.525 119.16 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.195 7.995 120.525 8.325 ;
        RECT 120.195 2.555 120.525 2.885 ;
        RECT 120.195 1.195 120.525 1.525 ;
        RECT 120.195 -0.165 120.525 0.165 ;
        RECT 120.195 -1.525 120.525 -1.195 ;
        RECT 120.2 -1.525 120.52 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 121.555 7.995 121.885 8.325 ;
        RECT 121.555 2.555 121.885 2.885 ;
        RECT 121.555 1.195 121.885 1.525 ;
        RECT 121.555 -0.165 121.885 0.165 ;
        RECT 121.555 -1.525 121.885 -1.195 ;
        RECT 121.56 -1.525 121.88 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.915 7.995 123.245 8.325 ;
        RECT 122.915 2.555 123.245 2.885 ;
        RECT 122.915 1.195 123.245 1.525 ;
        RECT 122.915 -0.165 123.245 0.165 ;
        RECT 122.915 -1.525 123.245 -1.195 ;
        RECT 122.92 -1.525 123.24 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.275 7.995 124.605 8.325 ;
        RECT 124.275 2.555 124.605 2.885 ;
        RECT 124.275 1.195 124.605 1.525 ;
        RECT 124.275 -0.165 124.605 0.165 ;
        RECT 124.275 -1.525 124.605 -1.195 ;
        RECT 124.28 -1.525 124.6 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.635 7.995 125.965 8.325 ;
        RECT 125.635 2.555 125.965 2.885 ;
        RECT 125.635 1.195 125.965 1.525 ;
        RECT 125.635 -0.165 125.965 0.165 ;
        RECT 125.635 -1.525 125.965 -1.195 ;
        RECT 125.64 -1.525 125.96 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.995 7.995 127.325 8.325 ;
        RECT 126.995 2.555 127.325 2.885 ;
        RECT 126.995 1.195 127.325 1.525 ;
        RECT 126.995 -0.165 127.325 0.165 ;
        RECT 126.995 -1.525 127.325 -1.195 ;
        RECT 127 -1.525 127.32 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.355 7.995 128.685 8.325 ;
        RECT 128.355 2.555 128.685 2.885 ;
        RECT 128.355 1.195 128.685 1.525 ;
        RECT 128.355 -0.165 128.685 0.165 ;
        RECT 128.355 -1.525 128.685 -1.195 ;
        RECT 128.36 -1.525 128.68 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.715 7.995 130.045 8.325 ;
        RECT 129.715 2.555 130.045 2.885 ;
        RECT 129.715 1.195 130.045 1.525 ;
        RECT 129.715 -0.165 130.045 0.165 ;
        RECT 129.715 -1.525 130.045 -1.195 ;
        RECT 129.72 -1.525 130.04 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.075 7.995 131.405 8.325 ;
        RECT 131.075 2.555 131.405 2.885 ;
        RECT 131.075 1.195 131.405 1.525 ;
        RECT 131.075 -0.165 131.405 0.165 ;
        RECT 131.075 -1.525 131.405 -1.195 ;
        RECT 131.08 -1.525 131.4 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.435 7.995 132.765 8.325 ;
        RECT 132.435 2.555 132.765 2.885 ;
        RECT 132.435 1.195 132.765 1.525 ;
        RECT 132.435 -0.165 132.765 0.165 ;
        RECT 132.435 -1.525 132.765 -1.195 ;
        RECT 132.44 -1.525 132.76 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.795 7.995 134.125 8.325 ;
        RECT 133.795 2.555 134.125 2.885 ;
        RECT 133.795 1.195 134.125 1.525 ;
        RECT 133.795 -0.165 134.125 0.165 ;
        RECT 133.795 -1.525 134.125 -1.195 ;
        RECT 133.8 -1.525 134.12 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.155 7.995 135.485 8.325 ;
        RECT 135.155 2.555 135.485 2.885 ;
        RECT 135.155 1.195 135.485 1.525 ;
        RECT 135.155 -0.165 135.485 0.165 ;
        RECT 135.155 -1.525 135.485 -1.195 ;
        RECT 135.16 -1.525 135.48 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 136.515 7.995 136.845 8.325 ;
        RECT 136.515 2.555 136.845 2.885 ;
        RECT 136.515 1.195 136.845 1.525 ;
        RECT 136.515 -0.165 136.845 0.165 ;
        RECT 136.515 -1.525 136.845 -1.195 ;
        RECT 136.52 -1.525 136.84 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.875 7.995 138.205 8.325 ;
        RECT 137.875 2.555 138.205 2.885 ;
        RECT 137.875 1.195 138.205 1.525 ;
        RECT 137.875 -0.165 138.205 0.165 ;
        RECT 137.875 -1.525 138.205 -1.195 ;
        RECT 137.88 -1.525 138.2 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.235 7.995 139.565 8.325 ;
        RECT 139.235 2.555 139.565 2.885 ;
        RECT 139.235 1.195 139.565 1.525 ;
        RECT 139.235 -0.165 139.565 0.165 ;
        RECT 139.235 -1.525 139.565 -1.195 ;
        RECT 139.24 -1.525 139.56 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.595 7.995 140.925 8.325 ;
        RECT 140.595 2.555 140.925 2.885 ;
        RECT 140.595 1.195 140.925 1.525 ;
        RECT 140.595 -0.165 140.925 0.165 ;
        RECT 140.595 -1.525 140.925 -1.195 ;
        RECT 140.6 -1.525 140.92 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.955 7.995 142.285 8.325 ;
        RECT 141.955 2.555 142.285 2.885 ;
        RECT 141.955 1.195 142.285 1.525 ;
        RECT 141.955 -0.165 142.285 0.165 ;
        RECT 141.955 -1.525 142.285 -1.195 ;
        RECT 141.96 -1.525 142.28 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.315 7.995 143.645 8.325 ;
        RECT 143.315 2.555 143.645 2.885 ;
        RECT 143.315 1.195 143.645 1.525 ;
        RECT 143.315 -0.165 143.645 0.165 ;
        RECT 143.315 -1.525 143.645 -1.195 ;
        RECT 143.32 -1.525 143.64 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 144.675 7.995 145.005 8.325 ;
        RECT 144.675 2.555 145.005 2.885 ;
        RECT 144.675 1.195 145.005 1.525 ;
        RECT 144.675 -0.165 145.005 0.165 ;
        RECT 144.675 -1.525 145.005 -1.195 ;
        RECT 144.68 -1.525 145 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.035 7.995 146.365 8.325 ;
        RECT 146.035 2.555 146.365 2.885 ;
        RECT 146.035 1.195 146.365 1.525 ;
        RECT 146.035 -0.165 146.365 0.165 ;
        RECT 146.035 -1.525 146.365 -1.195 ;
        RECT 146.04 -1.525 146.36 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.395 7.995 147.725 8.325 ;
        RECT 147.395 2.555 147.725 2.885 ;
        RECT 147.395 1.195 147.725 1.525 ;
        RECT 147.395 -0.165 147.725 0.165 ;
        RECT 147.395 -1.525 147.725 -1.195 ;
        RECT 147.4 -1.525 147.72 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.755 7.995 149.085 8.325 ;
        RECT 148.755 2.555 149.085 2.885 ;
        RECT 148.755 1.195 149.085 1.525 ;
        RECT 148.755 -0.165 149.085 0.165 ;
        RECT 148.755 -1.525 149.085 -1.195 ;
        RECT 148.76 -1.525 149.08 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.115 7.995 150.445 8.325 ;
        RECT 150.115 2.555 150.445 2.885 ;
        RECT 150.115 1.195 150.445 1.525 ;
        RECT 150.115 -0.165 150.445 0.165 ;
        RECT 150.115 -1.525 150.445 -1.195 ;
        RECT 150.12 -1.525 150.44 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 151.475 7.995 151.805 8.325 ;
        RECT 151.475 2.555 151.805 2.885 ;
        RECT 151.475 1.195 151.805 1.525 ;
        RECT 151.475 -0.165 151.805 0.165 ;
        RECT 151.475 -1.525 151.805 -1.195 ;
        RECT 151.48 -1.525 151.8 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.835 7.995 153.165 8.325 ;
        RECT 152.835 2.555 153.165 2.885 ;
        RECT 152.835 1.195 153.165 1.525 ;
        RECT 152.835 -0.165 153.165 0.165 ;
        RECT 152.835 -1.525 153.165 -1.195 ;
        RECT 152.84 -1.525 153.16 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.195 7.995 154.525 8.325 ;
        RECT 154.195 2.555 154.525 2.885 ;
        RECT 154.195 1.195 154.525 1.525 ;
        RECT 154.195 -0.165 154.525 0.165 ;
        RECT 154.195 -1.525 154.525 -1.195 ;
        RECT 154.2 -1.525 154.52 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.555 7.995 155.885 8.325 ;
        RECT 155.555 2.555 155.885 2.885 ;
        RECT 155.555 1.195 155.885 1.525 ;
        RECT 155.555 -0.165 155.885 0.165 ;
        RECT 155.555 -1.525 155.885 -1.195 ;
        RECT 155.56 -1.525 155.88 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.915 7.995 157.245 8.325 ;
        RECT 156.915 2.555 157.245 2.885 ;
        RECT 156.915 1.195 157.245 1.525 ;
        RECT 156.915 -0.165 157.245 0.165 ;
        RECT 156.915 -1.525 157.245 -1.195 ;
        RECT 156.92 -1.525 157.24 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.275 7.995 158.605 8.325 ;
        RECT 158.275 2.555 158.605 2.885 ;
        RECT 158.275 1.195 158.605 1.525 ;
        RECT 158.275 -0.165 158.605 0.165 ;
        RECT 158.275 -1.525 158.605 -1.195 ;
        RECT 158.28 -1.525 158.6 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.635 7.995 159.965 8.325 ;
        RECT 159.635 2.555 159.965 2.885 ;
        RECT 159.635 1.195 159.965 1.525 ;
        RECT 159.635 -0.165 159.965 0.165 ;
        RECT 159.635 -1.525 159.965 -1.195 ;
        RECT 159.64 -1.525 159.96 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.995 7.995 161.325 8.325 ;
        RECT 160.995 2.555 161.325 2.885 ;
        RECT 160.995 1.195 161.325 1.525 ;
        RECT 160.995 -0.165 161.325 0.165 ;
        RECT 160.995 -1.525 161.325 -1.195 ;
        RECT 161 -1.525 161.32 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 162.355 7.995 162.685 8.325 ;
        RECT 162.355 2.555 162.685 2.885 ;
        RECT 162.355 1.195 162.685 1.525 ;
        RECT 162.355 -0.165 162.685 0.165 ;
        RECT 162.355 -1.525 162.685 -1.195 ;
        RECT 162.36 -1.525 162.68 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.715 7.995 164.045 8.325 ;
        RECT 163.715 2.555 164.045 2.885 ;
        RECT 163.715 1.195 164.045 1.525 ;
        RECT 163.715 -0.165 164.045 0.165 ;
        RECT 163.715 -1.525 164.045 -1.195 ;
        RECT 163.72 -1.525 164.04 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.075 7.995 165.405 8.325 ;
        RECT 165.075 2.555 165.405 2.885 ;
        RECT 165.075 1.195 165.405 1.525 ;
        RECT 165.075 -0.165 165.405 0.165 ;
        RECT 165.075 -1.525 165.405 -1.195 ;
        RECT 165.08 -1.525 165.4 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.435 7.995 166.765 8.325 ;
        RECT 166.435 2.555 166.765 2.885 ;
        RECT 166.435 1.195 166.765 1.525 ;
        RECT 166.435 -0.165 166.765 0.165 ;
        RECT 166.435 -1.525 166.765 -1.195 ;
        RECT 166.44 -1.525 166.76 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.795 7.995 168.125 8.325 ;
        RECT 167.795 2.555 168.125 2.885 ;
        RECT 167.795 1.195 168.125 1.525 ;
        RECT 167.795 -0.165 168.125 0.165 ;
        RECT 167.795 -1.525 168.125 -1.195 ;
        RECT 167.8 -1.525 168.12 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.155 7.995 169.485 8.325 ;
        RECT 169.155 2.555 169.485 2.885 ;
        RECT 169.155 1.195 169.485 1.525 ;
        RECT 169.155 -0.165 169.485 0.165 ;
        RECT 169.155 -1.525 169.485 -1.195 ;
        RECT 169.16 -1.525 169.48 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.515 7.995 170.845 8.325 ;
        RECT 170.515 2.555 170.845 2.885 ;
        RECT 170.515 1.195 170.845 1.525 ;
        RECT 170.515 -0.165 170.845 0.165 ;
        RECT 170.515 -1.525 170.845 -1.195 ;
        RECT 170.52 -1.525 170.84 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.875 7.995 172.205 8.325 ;
        RECT 171.875 2.555 172.205 2.885 ;
        RECT 171.875 1.195 172.205 1.525 ;
        RECT 171.875 -0.165 172.205 0.165 ;
        RECT 171.875 -1.525 172.205 -1.195 ;
        RECT 171.88 -1.525 172.2 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.235 7.995 173.565 8.325 ;
        RECT 173.235 2.555 173.565 2.885 ;
        RECT 173.235 1.195 173.565 1.525 ;
        RECT 173.235 -0.165 173.565 0.165 ;
        RECT 173.235 -1.525 173.565 -1.195 ;
        RECT 173.24 -1.525 173.56 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 174.595 7.995 174.925 8.325 ;
        RECT 174.595 2.555 174.925 2.885 ;
        RECT 174.595 1.195 174.925 1.525 ;
        RECT 174.595 -0.165 174.925 0.165 ;
        RECT 174.595 -1.525 174.925 -1.195 ;
        RECT 174.6 -1.525 174.92 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.955 7.995 176.285 8.325 ;
        RECT 175.955 2.555 176.285 2.885 ;
        RECT 175.955 1.195 176.285 1.525 ;
        RECT 175.955 -0.165 176.285 0.165 ;
        RECT 175.955 -1.525 176.285 -1.195 ;
        RECT 175.96 -1.525 176.28 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.315 7.995 177.645 8.325 ;
        RECT 177.315 2.555 177.645 2.885 ;
        RECT 177.315 1.195 177.645 1.525 ;
        RECT 177.315 -0.165 177.645 0.165 ;
        RECT 177.315 -1.525 177.645 -1.195 ;
        RECT 177.32 -1.525 177.64 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 178.675 7.995 179.005 8.325 ;
        RECT 178.675 2.555 179.005 2.885 ;
        RECT 178.675 1.195 179.005 1.525 ;
        RECT 178.675 -0.165 179.005 0.165 ;
        RECT 178.675 -1.525 179.005 -1.195 ;
        RECT 178.68 -1.525 179 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.035 7.995 180.365 8.325 ;
        RECT 180.035 2.555 180.365 2.885 ;
        RECT 180.035 1.195 180.365 1.525 ;
        RECT 180.035 -0.165 180.365 0.165 ;
        RECT 180.035 -1.525 180.365 -1.195 ;
        RECT 180.04 -1.525 180.36 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 181.395 7.995 181.725 8.325 ;
        RECT 181.395 2.555 181.725 2.885 ;
        RECT 181.395 1.195 181.725 1.525 ;
        RECT 181.395 -0.165 181.725 0.165 ;
        RECT 181.395 -1.525 181.725 -1.195 ;
        RECT 181.4 -1.525 181.72 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.755 7.995 183.085 8.325 ;
        RECT 182.755 2.555 183.085 2.885 ;
        RECT 182.755 1.195 183.085 1.525 ;
        RECT 182.755 -0.165 183.085 0.165 ;
        RECT 182.755 -1.525 183.085 -1.195 ;
        RECT 182.76 -1.525 183.08 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.115 7.995 184.445 8.325 ;
        RECT 184.115 2.555 184.445 2.885 ;
        RECT 184.115 1.195 184.445 1.525 ;
        RECT 184.115 -0.165 184.445 0.165 ;
        RECT 184.115 -1.525 184.445 -1.195 ;
        RECT 184.12 -1.525 184.44 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 185.475 7.995 185.805 8.325 ;
        RECT 185.475 2.555 185.805 2.885 ;
        RECT 185.475 1.195 185.805 1.525 ;
        RECT 185.475 -0.165 185.805 0.165 ;
        RECT 185.475 -1.525 185.805 -1.195 ;
        RECT 185.48 -1.525 185.8 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.835 7.995 187.165 8.325 ;
        RECT 186.835 2.555 187.165 2.885 ;
        RECT 186.835 1.195 187.165 1.525 ;
        RECT 186.835 -0.165 187.165 0.165 ;
        RECT 186.835 -1.525 187.165 -1.195 ;
        RECT 186.84 -1.525 187.16 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.195 7.995 188.525 8.325 ;
        RECT 188.195 2.555 188.525 2.885 ;
        RECT 188.195 1.195 188.525 1.525 ;
        RECT 188.195 -0.165 188.525 0.165 ;
        RECT 188.195 -1.525 188.525 -1.195 ;
        RECT 188.2 -1.525 188.52 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.555 7.995 189.885 8.325 ;
        RECT 189.555 2.555 189.885 2.885 ;
        RECT 189.555 1.195 189.885 1.525 ;
        RECT 189.555 -0.165 189.885 0.165 ;
        RECT 189.555 -1.525 189.885 -1.195 ;
        RECT 189.56 -1.525 189.88 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.915 7.995 191.245 8.325 ;
        RECT 190.915 2.555 191.245 2.885 ;
        RECT 190.915 1.195 191.245 1.525 ;
        RECT 190.915 -0.165 191.245 0.165 ;
        RECT 190.915 -1.525 191.245 -1.195 ;
        RECT 190.92 -1.525 191.24 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.275 7.995 192.605 8.325 ;
        RECT 192.275 2.555 192.605 2.885 ;
        RECT 192.275 1.195 192.605 1.525 ;
        RECT 192.275 -0.165 192.605 0.165 ;
        RECT 192.275 -1.525 192.605 -1.195 ;
        RECT 192.28 -1.525 192.6 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 193.635 7.995 193.965 8.325 ;
        RECT 193.635 2.555 193.965 2.885 ;
        RECT 193.635 1.195 193.965 1.525 ;
        RECT 193.635 -0.165 193.965 0.165 ;
        RECT 193.635 -1.525 193.965 -1.195 ;
        RECT 193.64 -1.525 193.96 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.995 7.995 195.325 8.325 ;
        RECT 194.995 2.555 195.325 2.885 ;
        RECT 194.995 1.195 195.325 1.525 ;
        RECT 194.995 -0.165 195.325 0.165 ;
        RECT 194.995 -1.525 195.325 -1.195 ;
        RECT 195 -1.525 195.32 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 196.355 7.995 196.685 8.325 ;
        RECT 196.355 2.555 196.685 2.885 ;
        RECT 196.355 1.195 196.685 1.525 ;
        RECT 196.355 -0.165 196.685 0.165 ;
        RECT 196.355 -1.525 196.685 -1.195 ;
        RECT 196.36 -1.525 196.68 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.715 7.995 198.045 8.325 ;
        RECT 197.715 2.555 198.045 2.885 ;
        RECT 197.715 1.195 198.045 1.525 ;
        RECT 197.715 -0.165 198.045 0.165 ;
        RECT 197.715 -1.525 198.045 -1.195 ;
        RECT 197.72 -1.525 198.04 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.075 7.995 199.405 8.325 ;
        RECT 199.075 2.555 199.405 2.885 ;
        RECT 199.075 1.195 199.405 1.525 ;
        RECT 199.075 -0.165 199.405 0.165 ;
        RECT 199.075 -1.525 199.405 -1.195 ;
        RECT 199.08 -1.525 199.4 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 200.435 7.995 200.765 8.325 ;
        RECT 200.435 2.555 200.765 2.885 ;
        RECT 200.435 1.195 200.765 1.525 ;
        RECT 200.435 -0.165 200.765 0.165 ;
        RECT 200.435 -1.525 200.765 -1.195 ;
        RECT 200.44 -1.525 200.76 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.795 7.995 202.125 8.325 ;
        RECT 201.795 2.555 202.125 2.885 ;
        RECT 201.795 1.195 202.125 1.525 ;
        RECT 201.795 -0.165 202.125 0.165 ;
        RECT 201.795 -1.525 202.125 -1.195 ;
        RECT 201.8 -1.525 202.12 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.155 7.995 203.485 8.325 ;
        RECT 203.155 2.555 203.485 2.885 ;
        RECT 203.155 1.195 203.485 1.525 ;
        RECT 203.155 -0.165 203.485 0.165 ;
        RECT 203.155 -1.525 203.485 -1.195 ;
        RECT 203.16 -1.525 203.48 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 204.515 7.995 204.845 8.325 ;
        RECT 204.515 2.555 204.845 2.885 ;
        RECT 204.515 1.195 204.845 1.525 ;
        RECT 204.515 -0.165 204.845 0.165 ;
        RECT 204.515 -1.525 204.845 -1.195 ;
        RECT 204.52 -1.525 204.84 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.875 7.995 206.205 8.325 ;
        RECT 205.875 2.555 206.205 2.885 ;
        RECT 205.875 1.195 206.205 1.525 ;
        RECT 205.875 -0.165 206.205 0.165 ;
        RECT 205.875 -1.525 206.205 -1.195 ;
        RECT 205.88 -1.525 206.2 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.235 7.995 207.565 8.325 ;
        RECT 207.235 2.555 207.565 2.885 ;
        RECT 207.235 1.195 207.565 1.525 ;
        RECT 207.235 -0.165 207.565 0.165 ;
        RECT 207.235 -1.525 207.565 -1.195 ;
        RECT 207.24 -1.525 207.56 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 208.595 7.995 208.925 8.325 ;
        RECT 208.595 2.555 208.925 2.885 ;
        RECT 208.595 1.195 208.925 1.525 ;
        RECT 208.595 -0.165 208.925 0.165 ;
        RECT 208.595 -1.525 208.925 -1.195 ;
        RECT 208.6 -1.525 208.92 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.955 7.995 210.285 8.325 ;
        RECT 209.955 2.555 210.285 2.885 ;
        RECT 209.955 1.195 210.285 1.525 ;
        RECT 209.955 -0.165 210.285 0.165 ;
        RECT 209.955 -1.525 210.285 -1.195 ;
        RECT 209.96 -1.525 210.28 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 211.315 7.995 211.645 8.325 ;
        RECT 211.315 2.555 211.645 2.885 ;
        RECT 211.315 1.195 211.645 1.525 ;
        RECT 211.315 -0.165 211.645 0.165 ;
        RECT 211.315 -1.525 211.645 -1.195 ;
        RECT 211.32 -1.525 211.64 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 212.675 7.995 213.005 8.325 ;
        RECT 212.675 2.555 213.005 2.885 ;
        RECT 212.675 1.195 213.005 1.525 ;
        RECT 212.675 -0.165 213.005 0.165 ;
        RECT 212.675 -1.525 213.005 -1.195 ;
        RECT 212.68 -1.525 213 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.035 7.995 214.365 8.325 ;
        RECT 214.035 2.555 214.365 2.885 ;
        RECT 214.035 1.195 214.365 1.525 ;
        RECT 214.035 -0.165 214.365 0.165 ;
        RECT 214.035 -1.525 214.365 -1.195 ;
        RECT 214.04 -1.525 214.36 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 215.395 7.995 215.725 8.325 ;
        RECT 215.395 2.555 215.725 2.885 ;
        RECT 215.395 1.195 215.725 1.525 ;
        RECT 215.395 -0.165 215.725 0.165 ;
        RECT 215.395 -1.525 215.725 -1.195 ;
        RECT 215.4 -1.525 215.72 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.755 7.995 217.085 8.325 ;
        RECT 216.755 2.555 217.085 2.885 ;
        RECT 216.755 1.195 217.085 1.525 ;
        RECT 216.755 -0.165 217.085 0.165 ;
        RECT 216.755 -1.525 217.085 -1.195 ;
        RECT 216.76 -1.525 217.08 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.115 7.995 218.445 8.325 ;
        RECT 218.115 2.555 218.445 2.885 ;
        RECT 218.115 1.195 218.445 1.525 ;
        RECT 218.115 -0.165 218.445 0.165 ;
        RECT 218.115 -1.525 218.445 -1.195 ;
        RECT 218.12 -1.525 218.44 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 219.475 7.995 219.805 8.325 ;
        RECT 219.475 2.555 219.805 2.885 ;
        RECT 219.475 1.195 219.805 1.525 ;
        RECT 219.475 -0.165 219.805 0.165 ;
        RECT 219.475 -1.525 219.805 -1.195 ;
        RECT 219.48 -1.525 219.8 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.835 7.995 221.165 8.325 ;
        RECT 220.835 2.555 221.165 2.885 ;
        RECT 220.835 1.195 221.165 1.525 ;
        RECT 220.835 -0.165 221.165 0.165 ;
        RECT 220.835 -1.525 221.165 -1.195 ;
        RECT 220.84 -1.525 221.16 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.195 7.995 222.525 8.325 ;
        RECT 222.195 2.555 222.525 2.885 ;
        RECT 222.195 1.195 222.525 1.525 ;
        RECT 222.195 -0.165 222.525 0.165 ;
        RECT 222.195 -1.525 222.525 -1.195 ;
        RECT 222.2 -1.525 222.52 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 223.555 7.995 223.885 8.325 ;
        RECT 223.555 2.555 223.885 2.885 ;
        RECT 223.555 1.195 223.885 1.525 ;
        RECT 223.555 -0.165 223.885 0.165 ;
        RECT 223.555 -1.525 223.885 -1.195 ;
        RECT 223.56 -1.525 223.88 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 224.915 7.995 225.245 8.325 ;
        RECT 224.915 2.555 225.245 2.885 ;
        RECT 224.915 1.195 225.245 1.525 ;
        RECT 224.915 -0.165 225.245 0.165 ;
        RECT 224.915 -1.525 225.245 -1.195 ;
        RECT 224.92 -1.525 225.24 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.275 7.995 226.605 8.325 ;
        RECT 226.275 2.555 226.605 2.885 ;
        RECT 226.275 1.195 226.605 1.525 ;
        RECT 226.275 -0.165 226.605 0.165 ;
        RECT 226.275 -1.525 226.605 -1.195 ;
        RECT 226.28 -1.525 226.6 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 227.635 7.995 227.965 8.325 ;
        RECT 227.635 2.555 227.965 2.885 ;
        RECT 227.635 1.195 227.965 1.525 ;
        RECT 227.635 -0.165 227.965 0.165 ;
        RECT 227.635 -1.525 227.965 -1.195 ;
        RECT 227.64 -1.525 227.96 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.995 7.995 229.325 8.325 ;
        RECT 228.995 2.555 229.325 2.885 ;
        RECT 228.995 1.195 229.325 1.525 ;
        RECT 228.995 -0.165 229.325 0.165 ;
        RECT 228.995 -1.525 229.325 -1.195 ;
        RECT 229 -1.525 229.32 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 230.355 7.995 230.685 8.325 ;
        RECT 230.355 2.555 230.685 2.885 ;
        RECT 230.355 1.195 230.685 1.525 ;
        RECT 230.355 -0.165 230.685 0.165 ;
        RECT 230.355 -1.525 230.685 -1.195 ;
        RECT 230.36 -1.525 230.68 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 231.715 7.995 232.045 8.325 ;
        RECT 231.715 2.555 232.045 2.885 ;
        RECT 231.715 1.195 232.045 1.525 ;
        RECT 231.715 -0.165 232.045 0.165 ;
        RECT 231.715 -1.525 232.045 -1.195 ;
        RECT 231.72 -1.525 232.04 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.075 7.995 233.405 8.325 ;
        RECT 233.075 2.555 233.405 2.885 ;
        RECT 233.075 1.195 233.405 1.525 ;
        RECT 233.075 -0.165 233.405 0.165 ;
        RECT 233.075 -1.525 233.405 -1.195 ;
        RECT 233.08 -1.525 233.4 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 234.435 7.995 234.765 8.325 ;
        RECT 234.435 2.555 234.765 2.885 ;
        RECT 234.435 1.195 234.765 1.525 ;
        RECT 234.435 -0.165 234.765 0.165 ;
        RECT 234.435 -1.525 234.765 -1.195 ;
        RECT 234.44 -1.525 234.76 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 235.795 7.995 236.125 8.325 ;
        RECT 235.795 2.555 236.125 2.885 ;
        RECT 235.795 1.195 236.125 1.525 ;
        RECT 235.795 -0.165 236.125 0.165 ;
        RECT 235.795 -1.525 236.125 -1.195 ;
        RECT 235.8 -1.525 236.12 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 237.155 7.995 237.485 8.325 ;
        RECT 237.155 2.555 237.485 2.885 ;
        RECT 237.155 1.195 237.485 1.525 ;
        RECT 237.155 -0.165 237.485 0.165 ;
        RECT 237.155 -1.525 237.485 -1.195 ;
        RECT 237.16 -1.525 237.48 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 238.515 7.995 238.845 8.325 ;
        RECT 238.515 2.555 238.845 2.885 ;
        RECT 238.515 1.195 238.845 1.525 ;
        RECT 238.515 -0.165 238.845 0.165 ;
        RECT 238.515 -1.525 238.845 -1.195 ;
        RECT 238.52 -1.525 238.84 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.875 7.995 240.205 8.325 ;
        RECT 239.875 2.555 240.205 2.885 ;
        RECT 239.875 1.195 240.205 1.525 ;
        RECT 239.875 -0.165 240.205 0.165 ;
        RECT 239.875 -1.525 240.205 -1.195 ;
        RECT 239.88 -1.525 240.2 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 241.235 7.995 241.565 8.325 ;
        RECT 241.235 2.555 241.565 2.885 ;
        RECT 241.235 1.195 241.565 1.525 ;
        RECT 241.235 -0.165 241.565 0.165 ;
        RECT 241.235 -1.525 241.565 -1.195 ;
        RECT 241.24 -1.525 241.56 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 242.595 7.995 242.925 8.325 ;
        RECT 242.595 2.555 242.925 2.885 ;
        RECT 242.595 1.195 242.925 1.525 ;
        RECT 242.595 -0.165 242.925 0.165 ;
        RECT 242.595 -1.525 242.925 -1.195 ;
        RECT 242.6 -1.525 242.92 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 243.955 7.995 244.285 8.325 ;
        RECT 243.955 2.555 244.285 2.885 ;
        RECT 243.955 1.195 244.285 1.525 ;
        RECT 243.955 -0.165 244.285 0.165 ;
        RECT 243.955 -1.525 244.285 -1.195 ;
        RECT 243.96 -1.525 244.28 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 245.315 7.995 245.645 8.325 ;
        RECT 245.315 2.555 245.645 2.885 ;
        RECT 245.315 1.195 245.645 1.525 ;
        RECT 245.315 -0.165 245.645 0.165 ;
        RECT 245.315 -1.525 245.645 -1.195 ;
        RECT 245.32 -1.525 245.64 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 246.675 7.995 247.005 8.325 ;
        RECT 246.675 2.555 247.005 2.885 ;
        RECT 246.675 1.195 247.005 1.525 ;
        RECT 246.675 -0.165 247.005 0.165 ;
        RECT 246.675 -1.525 247.005 -1.195 ;
        RECT 246.68 -1.525 247 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.035 7.995 248.365 8.325 ;
        RECT 248.035 2.555 248.365 2.885 ;
        RECT 248.035 1.195 248.365 1.525 ;
        RECT 248.035 -0.165 248.365 0.165 ;
        RECT 248.035 -1.525 248.365 -1.195 ;
        RECT 248.04 -1.525 248.36 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 249.395 7.995 249.725 8.325 ;
        RECT 249.395 2.555 249.725 2.885 ;
        RECT 249.395 1.195 249.725 1.525 ;
        RECT 249.395 -0.165 249.725 0.165 ;
        RECT 249.395 -1.525 249.725 -1.195 ;
        RECT 249.4 -1.525 249.72 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.755 7.995 251.085 8.325 ;
        RECT 250.755 2.555 251.085 2.885 ;
        RECT 250.755 1.195 251.085 1.525 ;
        RECT 250.755 -0.165 251.085 0.165 ;
        RECT 250.755 -1.525 251.085 -1.195 ;
        RECT 250.76 -1.525 251.08 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.115 7.995 252.445 8.325 ;
        RECT 252.115 2.555 252.445 2.885 ;
        RECT 252.115 1.195 252.445 1.525 ;
        RECT 252.115 -0.165 252.445 0.165 ;
        RECT 252.115 -1.525 252.445 -1.195 ;
        RECT 252.12 -1.525 252.44 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 253.475 7.995 253.805 8.325 ;
        RECT 253.475 2.555 253.805 2.885 ;
        RECT 253.475 1.195 253.805 1.525 ;
        RECT 253.475 -0.165 253.805 0.165 ;
        RECT 253.475 -1.525 253.805 -1.195 ;
        RECT 253.48 -1.525 253.8 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 254.835 7.995 255.165 8.325 ;
        RECT 254.835 2.555 255.165 2.885 ;
        RECT 254.835 1.195 255.165 1.525 ;
        RECT 254.835 -0.165 255.165 0.165 ;
        RECT 254.835 -1.525 255.165 -1.195 ;
        RECT 254.84 -1.525 255.16 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 256.195 7.995 256.525 8.325 ;
        RECT 256.195 2.555 256.525 2.885 ;
        RECT 256.195 1.195 256.525 1.525 ;
        RECT 256.195 -0.165 256.525 0.165 ;
        RECT 256.195 -1.525 256.525 -1.195 ;
        RECT 256.2 -1.525 256.52 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 257.555 7.995 257.885 8.325 ;
        RECT 257.555 2.555 257.885 2.885 ;
        RECT 257.555 1.195 257.885 1.525 ;
        RECT 257.555 -0.165 257.885 0.165 ;
        RECT 257.555 -1.525 257.885 -1.195 ;
        RECT 257.56 -1.525 257.88 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.915 7.995 259.245 8.325 ;
        RECT 258.915 2.555 259.245 2.885 ;
        RECT 258.915 1.195 259.245 1.525 ;
        RECT 258.915 -0.165 259.245 0.165 ;
        RECT 258.915 -1.525 259.245 -1.195 ;
        RECT 258.92 -1.525 259.24 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.275 7.995 260.605 8.325 ;
        RECT 260.275 2.555 260.605 2.885 ;
        RECT 260.275 1.195 260.605 1.525 ;
        RECT 260.275 -0.165 260.605 0.165 ;
        RECT 260.275 -1.525 260.605 -1.195 ;
        RECT 260.28 -1.525 260.6 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 261.635 7.995 261.965 8.325 ;
        RECT 261.635 2.555 261.965 2.885 ;
        RECT 261.635 1.195 261.965 1.525 ;
        RECT 261.635 -0.165 261.965 0.165 ;
        RECT 261.635 -1.525 261.965 -1.195 ;
        RECT 261.64 -1.525 261.96 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.995 7.995 263.325 8.325 ;
        RECT 262.995 2.555 263.325 2.885 ;
        RECT 262.995 1.195 263.325 1.525 ;
        RECT 262.995 -0.165 263.325 0.165 ;
        RECT 262.995 -1.525 263.325 -1.195 ;
        RECT 263 -1.525 263.32 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 264.355 7.995 264.685 8.325 ;
        RECT 264.355 2.555 264.685 2.885 ;
        RECT 264.355 1.195 264.685 1.525 ;
        RECT 264.355 -0.165 264.685 0.165 ;
        RECT 264.355 -1.525 264.685 -1.195 ;
        RECT 264.36 -1.525 264.68 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 265.715 7.995 266.045 8.325 ;
        RECT 265.715 2.555 266.045 2.885 ;
        RECT 265.715 1.195 266.045 1.525 ;
        RECT 265.715 -0.165 266.045 0.165 ;
        RECT 265.715 -1.525 266.045 -1.195 ;
        RECT 265.72 -1.525 266.04 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 267.075 7.995 267.405 8.325 ;
        RECT 267.075 2.555 267.405 2.885 ;
        RECT 267.075 1.195 267.405 1.525 ;
        RECT 267.075 -0.165 267.405 0.165 ;
        RECT 267.075 -1.525 267.405 -1.195 ;
        RECT 267.08 -1.525 267.4 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 268.435 7.995 268.765 8.325 ;
        RECT 268.435 2.555 268.765 2.885 ;
        RECT 268.435 1.195 268.765 1.525 ;
        RECT 268.435 -0.165 268.765 0.165 ;
        RECT 268.435 -1.525 268.765 -1.195 ;
        RECT 268.44 -1.525 268.76 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.795 7.995 270.125 8.325 ;
        RECT 269.795 2.555 270.125 2.885 ;
        RECT 269.795 1.195 270.125 1.525 ;
        RECT 269.795 -0.165 270.125 0.165 ;
        RECT 269.795 -1.525 270.125 -1.195 ;
        RECT 269.8 -1.525 270.12 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.155 7.995 271.485 8.325 ;
        RECT 271.155 2.555 271.485 2.885 ;
        RECT 271.155 1.195 271.485 1.525 ;
        RECT 271.155 -0.165 271.485 0.165 ;
        RECT 271.155 -1.525 271.485 -1.195 ;
        RECT 271.16 -1.525 271.48 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 272.515 7.995 272.845 8.325 ;
        RECT 272.515 2.555 272.845 2.885 ;
        RECT 272.515 1.195 272.845 1.525 ;
        RECT 272.515 -0.165 272.845 0.165 ;
        RECT 272.515 -1.525 272.845 -1.195 ;
        RECT 272.52 -1.525 272.84 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.875 7.995 274.205 8.325 ;
        RECT 273.875 2.555 274.205 2.885 ;
        RECT 273.875 1.195 274.205 1.525 ;
        RECT 273.875 -0.165 274.205 0.165 ;
        RECT 273.875 -1.525 274.205 -1.195 ;
        RECT 273.88 -1.525 274.2 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.235 7.995 275.565 8.325 ;
        RECT 275.235 2.555 275.565 2.885 ;
        RECT 275.235 1.195 275.565 1.525 ;
        RECT 275.235 -0.165 275.565 0.165 ;
        RECT 275.235 -1.525 275.565 -1.195 ;
        RECT 275.24 -1.525 275.56 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 276.595 7.995 276.925 8.325 ;
        RECT 276.595 2.555 276.925 2.885 ;
        RECT 276.595 1.195 276.925 1.525 ;
        RECT 276.595 -0.165 276.925 0.165 ;
        RECT 276.595 -1.525 276.925 -1.195 ;
        RECT 276.6 -1.525 276.92 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 277.955 7.995 278.285 8.325 ;
        RECT 277.955 2.555 278.285 2.885 ;
        RECT 277.955 1.195 278.285 1.525 ;
        RECT 277.955 -0.165 278.285 0.165 ;
        RECT 277.955 -1.525 278.285 -1.195 ;
        RECT 277.96 -1.525 278.28 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.315 7.995 279.645 8.325 ;
        RECT 279.315 2.555 279.645 2.885 ;
        RECT 279.315 1.195 279.645 1.525 ;
        RECT 279.315 -0.165 279.645 0.165 ;
        RECT 279.315 -1.525 279.645 -1.195 ;
        RECT 279.32 -1.525 279.64 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 280.675 7.995 281.005 8.325 ;
        RECT 280.675 2.555 281.005 2.885 ;
        RECT 280.675 1.195 281.005 1.525 ;
        RECT 280.675 -0.165 281.005 0.165 ;
        RECT 280.675 -1.525 281.005 -1.195 ;
        RECT 280.68 -1.525 281 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.035 7.995 282.365 8.325 ;
        RECT 282.035 2.555 282.365 2.885 ;
        RECT 282.035 1.195 282.365 1.525 ;
        RECT 282.035 -0.165 282.365 0.165 ;
        RECT 282.035 -1.525 282.365 -1.195 ;
        RECT 282.04 -1.525 282.36 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 283.395 7.995 283.725 8.325 ;
        RECT 283.395 2.555 283.725 2.885 ;
        RECT 283.395 1.195 283.725 1.525 ;
        RECT 283.395 -0.165 283.725 0.165 ;
        RECT 283.395 -1.525 283.725 -1.195 ;
        RECT 283.4 -1.525 283.72 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 284.755 7.995 285.085 8.325 ;
        RECT 284.755 2.555 285.085 2.885 ;
        RECT 284.755 1.195 285.085 1.525 ;
        RECT 284.755 -0.165 285.085 0.165 ;
        RECT 284.755 -1.525 285.085 -1.195 ;
        RECT 284.76 -1.525 285.08 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.115 7.995 286.445 8.325 ;
        RECT 286.115 2.555 286.445 2.885 ;
        RECT 286.115 1.195 286.445 1.525 ;
        RECT 286.115 -0.165 286.445 0.165 ;
        RECT 286.115 -1.525 286.445 -1.195 ;
        RECT 286.12 -1.525 286.44 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 287.475 7.995 287.805 8.325 ;
        RECT 287.475 2.555 287.805 2.885 ;
        RECT 287.475 1.195 287.805 1.525 ;
        RECT 287.475 -0.165 287.805 0.165 ;
        RECT 287.475 -1.525 287.805 -1.195 ;
        RECT 287.48 -1.525 287.8 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.835 7.995 289.165 8.325 ;
        RECT 288.835 2.555 289.165 2.885 ;
        RECT 288.835 1.195 289.165 1.525 ;
        RECT 288.835 -0.165 289.165 0.165 ;
        RECT 288.835 -1.525 289.165 -1.195 ;
        RECT 288.84 -1.525 289.16 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.195 7.995 290.525 8.325 ;
        RECT 290.195 2.555 290.525 2.885 ;
        RECT 290.195 1.195 290.525 1.525 ;
        RECT 290.195 -0.165 290.525 0.165 ;
        RECT 290.195 -1.525 290.525 -1.195 ;
        RECT 290.2 -1.525 290.52 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 291.555 7.995 291.885 8.325 ;
        RECT 291.555 2.555 291.885 2.885 ;
        RECT 291.555 1.195 291.885 1.525 ;
        RECT 291.555 -0.165 291.885 0.165 ;
        RECT 291.555 -1.525 291.885 -1.195 ;
        RECT 291.56 -1.525 291.88 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.915 7.995 293.245 8.325 ;
        RECT 292.915 2.555 293.245 2.885 ;
        RECT 292.915 1.195 293.245 1.525 ;
        RECT 292.915 -0.165 293.245 0.165 ;
        RECT 292.915 -1.525 293.245 -1.195 ;
        RECT 292.92 -1.525 293.24 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.275 7.995 294.605 8.325 ;
        RECT 294.275 2.555 294.605 2.885 ;
        RECT 294.275 1.195 294.605 1.525 ;
        RECT 294.275 -0.165 294.605 0.165 ;
        RECT 294.275 -1.525 294.605 -1.195 ;
        RECT 294.28 -1.525 294.6 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 295.635 7.995 295.965 8.325 ;
        RECT 295.635 2.555 295.965 2.885 ;
        RECT 295.635 1.195 295.965 1.525 ;
        RECT 295.635 -0.165 295.965 0.165 ;
        RECT 295.635 -1.525 295.965 -1.195 ;
        RECT 295.64 -1.525 295.96 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 296.995 7.995 297.325 8.325 ;
        RECT 296.995 2.555 297.325 2.885 ;
        RECT 296.995 1.195 297.325 1.525 ;
        RECT 296.995 -0.165 297.325 0.165 ;
        RECT 296.995 -1.525 297.325 -1.195 ;
        RECT 297 -1.525 297.32 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 298.355 7.995 298.685 8.325 ;
        RECT 298.355 2.555 298.685 2.885 ;
        RECT 298.355 1.195 298.685 1.525 ;
        RECT 298.355 -0.165 298.685 0.165 ;
        RECT 298.355 -1.525 298.685 -1.195 ;
        RECT 298.36 -1.525 298.68 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 299.715 7.995 300.045 8.325 ;
        RECT 299.715 2.555 300.045 2.885 ;
        RECT 299.715 1.195 300.045 1.525 ;
        RECT 299.715 -0.165 300.045 0.165 ;
        RECT 299.715 -1.525 300.045 -1.195 ;
        RECT 299.72 -1.525 300.04 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.075 7.995 301.405 8.325 ;
        RECT 301.075 2.555 301.405 2.885 ;
        RECT 301.075 1.195 301.405 1.525 ;
        RECT 301.075 -0.165 301.405 0.165 ;
        RECT 301.075 -1.525 301.405 -1.195 ;
        RECT 301.08 -1.525 301.4 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 302.435 7.995 302.765 8.325 ;
        RECT 302.435 2.555 302.765 2.885 ;
        RECT 302.435 1.195 302.765 1.525 ;
        RECT 302.435 -0.165 302.765 0.165 ;
        RECT 302.435 -1.525 302.765 -1.195 ;
        RECT 302.44 -1.525 302.76 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.795 7.995 304.125 8.325 ;
        RECT 303.795 2.555 304.125 2.885 ;
        RECT 303.795 1.195 304.125 1.525 ;
        RECT 303.795 -0.165 304.125 0.165 ;
        RECT 303.795 -1.525 304.125 -1.195 ;
        RECT 303.8 -1.525 304.12 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.155 7.995 305.485 8.325 ;
        RECT 305.155 2.555 305.485 2.885 ;
        RECT 305.155 1.195 305.485 1.525 ;
        RECT 305.155 -0.165 305.485 0.165 ;
        RECT 305.155 -1.525 305.485 -1.195 ;
        RECT 305.16 -1.525 305.48 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 306.515 7.995 306.845 8.325 ;
        RECT 306.515 2.555 306.845 2.885 ;
        RECT 306.515 1.195 306.845 1.525 ;
        RECT 306.515 -0.165 306.845 0.165 ;
        RECT 306.515 -1.525 306.845 -1.195 ;
        RECT 306.52 -1.525 306.84 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.875 7.995 308.205 8.325 ;
        RECT 307.875 2.555 308.205 2.885 ;
        RECT 307.875 1.195 308.205 1.525 ;
        RECT 307.875 -0.165 308.205 0.165 ;
        RECT 307.875 -1.525 308.205 -1.195 ;
        RECT 307.88 -1.525 308.2 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.235 7.995 309.565 8.325 ;
        RECT 309.235 2.555 309.565 2.885 ;
        RECT 309.235 1.195 309.565 1.525 ;
        RECT 309.235 -0.165 309.565 0.165 ;
        RECT 309.235 -1.525 309.565 -1.195 ;
        RECT 309.24 -1.525 309.56 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 310.595 7.995 310.925 8.325 ;
        RECT 310.595 2.555 310.925 2.885 ;
        RECT 310.595 1.195 310.925 1.525 ;
        RECT 310.595 -0.165 310.925 0.165 ;
        RECT 310.595 -1.525 310.925 -1.195 ;
        RECT 310.6 -1.525 310.92 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 311.955 7.995 312.285 8.325 ;
        RECT 311.955 2.555 312.285 2.885 ;
        RECT 311.955 1.195 312.285 1.525 ;
        RECT 311.955 -0.165 312.285 0.165 ;
        RECT 311.955 -1.525 312.285 -1.195 ;
        RECT 311.96 -1.525 312.28 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.315 7.995 313.645 8.325 ;
        RECT 313.315 2.555 313.645 2.885 ;
        RECT 313.315 1.195 313.645 1.525 ;
        RECT 313.315 -0.165 313.645 0.165 ;
        RECT 313.315 -1.525 313.645 -1.195 ;
        RECT 313.32 -1.525 313.64 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 314.675 7.995 315.005 8.325 ;
        RECT 314.675 2.555 315.005 2.885 ;
        RECT 314.675 1.195 315.005 1.525 ;
        RECT 314.675 -0.165 315.005 0.165 ;
        RECT 314.675 -1.525 315.005 -1.195 ;
        RECT 314.68 -1.525 315 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 316.035 7.995 316.365 8.325 ;
        RECT 316.035 2.555 316.365 2.885 ;
        RECT 316.035 1.195 316.365 1.525 ;
        RECT 316.035 -0.165 316.365 0.165 ;
        RECT 316.035 -1.525 316.365 -1.195 ;
        RECT 316.04 -1.525 316.36 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 317.395 7.995 317.725 8.325 ;
        RECT 317.395 2.555 317.725 2.885 ;
        RECT 317.395 1.195 317.725 1.525 ;
        RECT 317.395 -0.165 317.725 0.165 ;
        RECT 317.395 -1.525 317.725 -1.195 ;
        RECT 317.4 -1.525 317.72 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.755 -0.165 319.085 0.165 ;
        RECT 318.755 -1.525 319.085 -1.195 ;
        RECT 318.76 -1.525 319.08 9 ;
        RECT 318.755 7.995 319.085 8.325 ;
        RECT 318.755 2.555 319.085 2.885 ;
        RECT 318.755 1.195 319.085 1.525 ;
    END
    PORT
      LAYER met3 ;
        RECT -2.205 7.995 -1.875 8.325 ;
        RECT -2.205 6.635 -1.875 6.965 ;
        RECT -2.205 5.275 -1.875 5.605 ;
        RECT -2.205 3.915 -1.875 4.245 ;
        RECT -2.205 2.555 -1.875 2.885 ;
        RECT -2.205 1.195 -1.875 1.525 ;
        RECT -2.205 -0.165 -1.875 0.165 ;
        RECT -2.205 -1.525 -1.875 -1.195 ;
        RECT -2.2 -1.525 -1.88 9 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.845 7.995 -0.515 8.325 ;
        RECT -0.845 6.635 -0.515 6.965 ;
        RECT -0.845 5.275 -0.515 5.605 ;
        RECT -0.845 3.915 -0.515 4.245 ;
        RECT -0.845 2.555 -0.515 2.885 ;
        RECT -0.845 1.195 -0.515 1.525 ;
        RECT -0.845 -0.165 -0.515 0.165 ;
        RECT -0.845 -1.525 -0.515 -1.195 ;
        RECT -0.84 -1.525 -0.52 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.515 7.995 0.845 8.325 ;
        RECT 0.515 5.275 0.845 5.605 ;
        RECT 0.515 3.915 0.845 4.245 ;
        RECT 0.515 2.555 0.845 2.885 ;
        RECT 0.515 1.195 0.845 1.525 ;
        RECT 0.515 -0.165 0.845 0.165 ;
        RECT 0.515 -1.525 0.845 -1.195 ;
        RECT 0.52 -1.525 0.84 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.875 7.995 2.205 8.325 ;
        RECT 1.875 5.275 2.205 5.605 ;
        RECT 1.875 2.555 2.205 2.885 ;
        RECT 1.875 1.195 2.205 1.525 ;
        RECT 1.875 -0.165 2.205 0.165 ;
        RECT 1.875 -1.525 2.205 -1.195 ;
        RECT 1.88 -1.525 2.2 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.235 7.995 3.565 8.325 ;
        RECT 3.235 5.275 3.565 5.605 ;
        RECT 3.235 2.555 3.565 2.885 ;
        RECT 3.235 1.195 3.565 1.525 ;
        RECT 3.235 -0.165 3.565 0.165 ;
        RECT 3.235 -1.525 3.565 -1.195 ;
        RECT 3.24 -1.525 3.56 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.595 7.995 4.925 8.325 ;
        RECT 4.595 2.555 4.925 2.885 ;
        RECT 4.595 1.195 4.925 1.525 ;
        RECT 4.595 -0.165 4.925 0.165 ;
        RECT 4.595 -1.525 4.925 -1.195 ;
        RECT 4.6 -1.525 4.92 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.955 7.995 6.285 8.325 ;
        RECT 5.955 2.555 6.285 2.885 ;
        RECT 5.955 1.195 6.285 1.525 ;
        RECT 5.955 -0.165 6.285 0.165 ;
        RECT 5.955 -1.525 6.285 -1.195 ;
        RECT 5.96 -1.525 6.28 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.315 7.995 7.645 8.325 ;
        RECT 7.315 2.555 7.645 2.885 ;
        RECT 7.315 1.195 7.645 1.525 ;
        RECT 7.315 -0.165 7.645 0.165 ;
        RECT 7.315 -1.525 7.645 -1.195 ;
        RECT 7.32 -1.525 7.64 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.675 7.995 9.005 8.325 ;
        RECT 8.675 2.555 9.005 2.885 ;
        RECT 8.675 1.195 9.005 1.525 ;
        RECT 8.675 -0.165 9.005 0.165 ;
        RECT 8.675 -1.525 9.005 -1.195 ;
        RECT 8.68 -1.525 9 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.035 7.995 10.365 8.325 ;
        RECT 10.035 2.555 10.365 2.885 ;
        RECT 10.035 1.195 10.365 1.525 ;
        RECT 10.035 -0.165 10.365 0.165 ;
        RECT 10.035 -1.525 10.365 -1.195 ;
        RECT 10.04 -1.525 10.36 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.395 7.995 11.725 8.325 ;
        RECT 11.395 2.555 11.725 2.885 ;
        RECT 11.395 1.195 11.725 1.525 ;
        RECT 11.395 -0.165 11.725 0.165 ;
        RECT 11.395 -1.525 11.725 -1.195 ;
        RECT 11.4 -1.525 11.72 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.755 7.995 13.085 8.325 ;
        RECT 12.755 2.555 13.085 2.885 ;
        RECT 12.755 1.195 13.085 1.525 ;
        RECT 12.755 -0.165 13.085 0.165 ;
        RECT 12.755 -1.525 13.085 -1.195 ;
        RECT 12.76 -1.525 13.08 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.115 7.995 14.445 8.325 ;
        RECT 14.115 2.555 14.445 2.885 ;
        RECT 14.115 1.195 14.445 1.525 ;
        RECT 14.115 -0.165 14.445 0.165 ;
        RECT 14.115 -1.525 14.445 -1.195 ;
        RECT 14.12 -1.525 14.44 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.475 7.995 15.805 8.325 ;
        RECT 15.475 2.555 15.805 2.885 ;
        RECT 15.475 1.195 15.805 1.525 ;
        RECT 15.475 -0.165 15.805 0.165 ;
        RECT 15.475 -1.525 15.805 -1.195 ;
        RECT 15.48 -1.525 15.8 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.835 7.995 17.165 8.325 ;
        RECT 16.835 2.555 17.165 2.885 ;
        RECT 16.835 1.195 17.165 1.525 ;
        RECT 16.835 -0.165 17.165 0.165 ;
        RECT 16.835 -1.525 17.165 -1.195 ;
        RECT 16.84 -1.525 17.16 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.195 7.995 18.525 8.325 ;
        RECT 18.195 2.555 18.525 2.885 ;
        RECT 18.195 1.195 18.525 1.525 ;
        RECT 18.195 -0.165 18.525 0.165 ;
        RECT 18.195 -1.525 18.525 -1.195 ;
        RECT 18.2 -1.525 18.52 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.555 7.995 19.885 8.325 ;
        RECT 19.555 2.555 19.885 2.885 ;
        RECT 19.555 1.195 19.885 1.525 ;
        RECT 19.555 -0.165 19.885 0.165 ;
        RECT 19.555 -1.525 19.885 -1.195 ;
        RECT 19.56 -1.525 19.88 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.915 7.995 21.245 8.325 ;
        RECT 20.915 2.555 21.245 2.885 ;
        RECT 20.915 1.195 21.245 1.525 ;
        RECT 20.915 -0.165 21.245 0.165 ;
        RECT 20.915 -1.525 21.245 -1.195 ;
        RECT 20.92 -1.525 21.24 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.275 7.995 22.605 8.325 ;
        RECT 22.275 2.555 22.605 2.885 ;
        RECT 22.275 1.195 22.605 1.525 ;
        RECT 22.275 -0.165 22.605 0.165 ;
        RECT 22.275 -1.525 22.605 -1.195 ;
        RECT 22.28 -1.525 22.6 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.635 7.995 23.965 8.325 ;
        RECT 23.635 2.555 23.965 2.885 ;
        RECT 23.635 1.195 23.965 1.525 ;
        RECT 23.635 -0.165 23.965 0.165 ;
        RECT 23.635 -1.525 23.965 -1.195 ;
        RECT 23.64 -1.525 23.96 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.995 7.995 25.325 8.325 ;
        RECT 24.995 2.555 25.325 2.885 ;
        RECT 24.995 1.195 25.325 1.525 ;
        RECT 24.995 -0.165 25.325 0.165 ;
        RECT 24.995 -1.525 25.325 -1.195 ;
        RECT 25 -1.525 25.32 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.355 7.995 26.685 8.325 ;
        RECT 26.355 2.555 26.685 2.885 ;
        RECT 26.355 1.195 26.685 1.525 ;
        RECT 26.355 -0.165 26.685 0.165 ;
        RECT 26.355 -1.525 26.685 -1.195 ;
        RECT 26.36 -1.525 26.68 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.715 7.995 28.045 8.325 ;
        RECT 27.715 2.555 28.045 2.885 ;
        RECT 27.715 1.195 28.045 1.525 ;
        RECT 27.715 -0.165 28.045 0.165 ;
        RECT 27.715 -1.525 28.045 -1.195 ;
        RECT 27.72 -1.525 28.04 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.075 7.995 29.405 8.325 ;
        RECT 29.075 2.555 29.405 2.885 ;
        RECT 29.075 1.195 29.405 1.525 ;
        RECT 29.075 -0.165 29.405 0.165 ;
        RECT 29.075 -1.525 29.405 -1.195 ;
        RECT 29.08 -1.525 29.4 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.435 7.995 30.765 8.325 ;
        RECT 30.435 2.555 30.765 2.885 ;
        RECT 30.435 1.195 30.765 1.525 ;
        RECT 30.435 -0.165 30.765 0.165 ;
        RECT 30.435 -1.525 30.765 -1.195 ;
        RECT 30.44 -1.525 30.76 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.795 7.995 32.125 8.325 ;
        RECT 31.795 2.555 32.125 2.885 ;
        RECT 31.795 1.195 32.125 1.525 ;
        RECT 31.795 -0.165 32.125 0.165 ;
        RECT 31.795 -1.525 32.125 -1.195 ;
        RECT 31.8 -1.525 32.12 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.155 7.995 33.485 8.325 ;
        RECT 33.155 2.555 33.485 2.885 ;
        RECT 33.155 1.195 33.485 1.525 ;
        RECT 33.155 -0.165 33.485 0.165 ;
        RECT 33.155 -1.525 33.485 -1.195 ;
        RECT 33.16 -1.525 33.48 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.515 7.995 34.845 8.325 ;
        RECT 34.515 2.555 34.845 2.885 ;
        RECT 34.515 1.195 34.845 1.525 ;
        RECT 34.515 -0.165 34.845 0.165 ;
        RECT 34.515 -1.525 34.845 -1.195 ;
        RECT 34.52 -1.525 34.84 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.875 7.995 36.205 8.325 ;
        RECT 35.875 2.555 36.205 2.885 ;
        RECT 35.875 1.195 36.205 1.525 ;
        RECT 35.875 -0.165 36.205 0.165 ;
        RECT 35.875 -1.525 36.205 -1.195 ;
        RECT 35.88 -1.525 36.2 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.235 7.995 37.565 8.325 ;
        RECT 37.235 2.555 37.565 2.885 ;
        RECT 37.235 1.195 37.565 1.525 ;
        RECT 37.235 -0.165 37.565 0.165 ;
        RECT 37.235 -1.525 37.565 -1.195 ;
        RECT 37.24 -1.525 37.56 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.595 7.995 38.925 8.325 ;
        RECT 38.595 2.555 38.925 2.885 ;
        RECT 38.595 1.195 38.925 1.525 ;
        RECT 38.595 -0.165 38.925 0.165 ;
        RECT 38.595 -1.525 38.925 -1.195 ;
        RECT 38.6 -1.525 38.92 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.955 7.995 40.285 8.325 ;
        RECT 39.955 2.555 40.285 2.885 ;
        RECT 39.955 1.195 40.285 1.525 ;
        RECT 39.955 -0.165 40.285 0.165 ;
        RECT 39.955 -1.525 40.285 -1.195 ;
        RECT 39.96 -1.525 40.28 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.315 7.995 41.645 8.325 ;
        RECT 41.315 2.555 41.645 2.885 ;
        RECT 41.315 1.195 41.645 1.525 ;
        RECT 41.315 -0.165 41.645 0.165 ;
        RECT 41.315 -1.525 41.645 -1.195 ;
        RECT 41.32 -1.525 41.64 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.675 7.995 43.005 8.325 ;
        RECT 42.675 2.555 43.005 2.885 ;
        RECT 42.675 1.195 43.005 1.525 ;
        RECT 42.675 -0.165 43.005 0.165 ;
        RECT 42.675 -1.525 43.005 -1.195 ;
        RECT 42.68 -1.525 43 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.035 7.995 44.365 8.325 ;
        RECT 44.035 2.555 44.365 2.885 ;
        RECT 44.035 1.195 44.365 1.525 ;
        RECT 44.035 -0.165 44.365 0.165 ;
        RECT 44.035 -1.525 44.365 -1.195 ;
        RECT 44.04 -1.525 44.36 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.395 7.995 45.725 8.325 ;
        RECT 45.395 2.555 45.725 2.885 ;
        RECT 45.395 1.195 45.725 1.525 ;
        RECT 45.395 -0.165 45.725 0.165 ;
        RECT 45.395 -1.525 45.725 -1.195 ;
        RECT 45.4 -1.525 45.72 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.755 7.995 47.085 8.325 ;
        RECT 46.755 2.555 47.085 2.885 ;
        RECT 46.755 1.195 47.085 1.525 ;
        RECT 46.755 -0.165 47.085 0.165 ;
        RECT 46.755 -1.525 47.085 -1.195 ;
        RECT 46.76 -1.525 47.08 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.115 7.995 48.445 8.325 ;
        RECT 48.115 2.555 48.445 2.885 ;
        RECT 48.115 1.195 48.445 1.525 ;
        RECT 48.115 -0.165 48.445 0.165 ;
        RECT 48.115 -1.525 48.445 -1.195 ;
        RECT 48.12 -1.525 48.44 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.475 7.995 49.805 8.325 ;
        RECT 49.475 2.555 49.805 2.885 ;
        RECT 49.475 1.195 49.805 1.525 ;
        RECT 49.475 -0.165 49.805 0.165 ;
        RECT 49.475 -1.525 49.805 -1.195 ;
        RECT 49.48 -1.525 49.8 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.835 7.995 51.165 8.325 ;
        RECT 50.835 2.555 51.165 2.885 ;
        RECT 50.835 1.195 51.165 1.525 ;
        RECT 50.835 -0.165 51.165 0.165 ;
        RECT 50.835 -1.525 51.165 -1.195 ;
        RECT 50.84 -1.525 51.16 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.195 7.995 52.525 8.325 ;
        RECT 52.195 2.555 52.525 2.885 ;
        RECT 52.195 1.195 52.525 1.525 ;
        RECT 52.195 -0.165 52.525 0.165 ;
        RECT 52.195 -1.525 52.525 -1.195 ;
        RECT 52.2 -1.525 52.52 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.555 7.995 53.885 8.325 ;
        RECT 53.555 2.555 53.885 2.885 ;
        RECT 53.555 1.195 53.885 1.525 ;
        RECT 53.555 -0.165 53.885 0.165 ;
        RECT 53.555 -1.525 53.885 -1.195 ;
        RECT 53.56 -1.525 53.88 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.915 7.995 55.245 8.325 ;
        RECT 54.915 2.555 55.245 2.885 ;
        RECT 54.915 1.195 55.245 1.525 ;
        RECT 54.915 -0.165 55.245 0.165 ;
        RECT 54.915 -1.525 55.245 -1.195 ;
        RECT 54.92 -1.525 55.24 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.275 7.995 56.605 8.325 ;
        RECT 56.275 2.555 56.605 2.885 ;
        RECT 56.275 1.195 56.605 1.525 ;
        RECT 56.275 -0.165 56.605 0.165 ;
        RECT 56.275 -1.525 56.605 -1.195 ;
        RECT 56.28 -1.525 56.6 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.635 7.995 57.965 8.325 ;
        RECT 57.635 2.555 57.965 2.885 ;
        RECT 57.635 1.195 57.965 1.525 ;
        RECT 57.635 -0.165 57.965 0.165 ;
        RECT 57.635 -1.525 57.965 -1.195 ;
        RECT 57.64 -1.525 57.96 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.995 7.995 59.325 8.325 ;
        RECT 58.995 2.555 59.325 2.885 ;
        RECT 58.995 1.195 59.325 1.525 ;
        RECT 58.995 -0.165 59.325 0.165 ;
        RECT 58.995 -1.525 59.325 -1.195 ;
        RECT 59 -1.525 59.32 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.355 7.995 60.685 8.325 ;
        RECT 60.355 2.555 60.685 2.885 ;
        RECT 60.355 1.195 60.685 1.525 ;
        RECT 60.355 -0.165 60.685 0.165 ;
        RECT 60.355 -1.525 60.685 -1.195 ;
        RECT 60.36 -1.525 60.68 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.715 7.995 62.045 8.325 ;
        RECT 61.715 2.555 62.045 2.885 ;
        RECT 61.715 1.195 62.045 1.525 ;
        RECT 61.715 -0.165 62.045 0.165 ;
        RECT 61.715 -1.525 62.045 -1.195 ;
        RECT 61.72 -1.525 62.04 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.075 7.995 63.405 8.325 ;
        RECT 63.075 2.555 63.405 2.885 ;
        RECT 63.075 1.195 63.405 1.525 ;
        RECT 63.075 -0.165 63.405 0.165 ;
        RECT 63.075 -1.525 63.405 -1.195 ;
        RECT 63.08 -1.525 63.4 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.435 7.995 64.765 8.325 ;
        RECT 64.435 2.555 64.765 2.885 ;
        RECT 64.435 1.195 64.765 1.525 ;
        RECT 64.435 -0.165 64.765 0.165 ;
        RECT 64.435 -1.525 64.765 -1.195 ;
        RECT 64.44 -1.525 64.76 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.795 7.995 66.125 8.325 ;
        RECT 65.795 2.555 66.125 2.885 ;
        RECT 65.795 1.195 66.125 1.525 ;
        RECT 65.795 -0.165 66.125 0.165 ;
        RECT 65.795 -1.525 66.125 -1.195 ;
        RECT 65.8 -1.525 66.12 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.155 7.995 67.485 8.325 ;
        RECT 67.155 2.555 67.485 2.885 ;
        RECT 67.155 1.195 67.485 1.525 ;
        RECT 67.155 -0.165 67.485 0.165 ;
        RECT 67.155 -1.525 67.485 -1.195 ;
        RECT 67.16 -1.525 67.48 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.515 7.995 68.845 8.325 ;
        RECT 68.515 2.555 68.845 2.885 ;
        RECT 68.515 1.195 68.845 1.525 ;
        RECT 68.515 -0.165 68.845 0.165 ;
        RECT 68.515 -1.525 68.845 -1.195 ;
        RECT 68.52 -1.525 68.84 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.875 7.995 70.205 8.325 ;
        RECT 69.875 2.555 70.205 2.885 ;
        RECT 69.875 1.195 70.205 1.525 ;
        RECT 69.875 -0.165 70.205 0.165 ;
        RECT 69.875 -1.525 70.205 -1.195 ;
        RECT 69.88 -1.525 70.2 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.235 7.995 71.565 8.325 ;
        RECT 71.235 2.555 71.565 2.885 ;
        RECT 71.235 1.195 71.565 1.525 ;
        RECT 71.235 -0.165 71.565 0.165 ;
        RECT 71.235 -1.525 71.565 -1.195 ;
        RECT 71.24 -1.525 71.56 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.595 7.995 72.925 8.325 ;
        RECT 72.595 2.555 72.925 2.885 ;
        RECT 72.595 1.195 72.925 1.525 ;
        RECT 72.595 -0.165 72.925 0.165 ;
        RECT 72.595 -1.525 72.925 -1.195 ;
        RECT 72.6 -1.525 72.92 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 7.995 74.285 8.325 ;
        RECT 73.955 2.555 74.285 2.885 ;
        RECT 73.955 1.195 74.285 1.525 ;
        RECT 73.955 -0.165 74.285 0.165 ;
        RECT 73.955 -1.525 74.285 -1.195 ;
        RECT 73.96 -1.525 74.28 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.315 7.995 75.645 8.325 ;
        RECT 75.315 2.555 75.645 2.885 ;
        RECT 75.315 1.195 75.645 1.525 ;
        RECT 75.315 -0.165 75.645 0.165 ;
        RECT 75.315 -1.525 75.645 -1.195 ;
        RECT 75.32 -1.525 75.64 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 76.675 7.995 77.005 8.325 ;
        RECT 76.675 2.555 77.005 2.885 ;
        RECT 76.675 1.195 77.005 1.525 ;
        RECT 76.675 -0.165 77.005 0.165 ;
        RECT 76.675 -1.525 77.005 -1.195 ;
        RECT 76.68 -1.525 77 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.035 7.995 78.365 8.325 ;
        RECT 78.035 2.555 78.365 2.885 ;
        RECT 78.035 1.195 78.365 1.525 ;
        RECT 78.035 -0.165 78.365 0.165 ;
        RECT 78.035 -1.525 78.365 -1.195 ;
        RECT 78.04 -1.525 78.36 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 79.395 7.995 79.725 8.325 ;
        RECT 79.395 2.555 79.725 2.885 ;
        RECT 79.395 1.195 79.725 1.525 ;
        RECT 79.395 -0.165 79.725 0.165 ;
        RECT 79.395 -1.525 79.725 -1.195 ;
        RECT 79.4 -1.525 79.72 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.755 7.995 81.085 8.325 ;
        RECT 80.755 2.555 81.085 2.885 ;
        RECT 80.755 1.195 81.085 1.525 ;
        RECT 80.755 -0.165 81.085 0.165 ;
        RECT 80.755 -1.525 81.085 -1.195 ;
        RECT 80.76 -1.525 81.08 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.115 7.995 82.445 8.325 ;
        RECT 82.115 2.555 82.445 2.885 ;
        RECT 82.115 1.195 82.445 1.525 ;
        RECT 82.115 -0.165 82.445 0.165 ;
        RECT 82.115 -1.525 82.445 -1.195 ;
        RECT 82.12 -1.525 82.44 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 83.475 7.995 83.805 8.325 ;
        RECT 83.475 2.555 83.805 2.885 ;
        RECT 83.475 1.195 83.805 1.525 ;
        RECT 83.475 -0.165 83.805 0.165 ;
        RECT 83.475 -1.525 83.805 -1.195 ;
        RECT 83.48 -1.525 83.8 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.835 7.995 85.165 8.325 ;
        RECT 84.835 2.555 85.165 2.885 ;
        RECT 84.835 1.195 85.165 1.525 ;
        RECT 84.835 -0.165 85.165 0.165 ;
        RECT 84.835 -1.525 85.165 -1.195 ;
        RECT 84.84 -1.525 85.16 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.195 7.995 86.525 8.325 ;
        RECT 86.195 2.555 86.525 2.885 ;
        RECT 86.195 1.195 86.525 1.525 ;
        RECT 86.195 -0.165 86.525 0.165 ;
        RECT 86.195 -1.525 86.525 -1.195 ;
        RECT 86.2 -1.525 86.52 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.555 7.995 87.885 8.325 ;
        RECT 87.555 2.555 87.885 2.885 ;
        RECT 87.555 1.195 87.885 1.525 ;
        RECT 87.555 -0.165 87.885 0.165 ;
        RECT 87.555 -1.525 87.885 -1.195 ;
        RECT 87.56 -1.525 87.88 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.915 7.995 89.245 8.325 ;
        RECT 88.915 2.555 89.245 2.885 ;
        RECT 88.915 1.195 89.245 1.525 ;
        RECT 88.915 -0.165 89.245 0.165 ;
        RECT 88.915 -1.525 89.245 -1.195 ;
        RECT 88.92 -1.525 89.24 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.275 7.995 90.605 8.325 ;
        RECT 90.275 2.555 90.605 2.885 ;
        RECT 90.275 1.195 90.605 1.525 ;
        RECT 90.275 -0.165 90.605 0.165 ;
        RECT 90.275 -1.525 90.605 -1.195 ;
        RECT 90.28 -1.525 90.6 9 ;
    END
    PORT
      LAYER met3 ;
        RECT 91.635 2.555 91.965 2.885 ;
        RECT 91.635 1.195 91.965 1.525 ;
        RECT 91.635 -0.165 91.965 0.165 ;
        RECT 91.635 -1.525 91.965 -1.195 ;
        RECT 91.64 -1.525 91.96 9 ;
        RECT 91.635 7.995 91.965 8.325 ;
    END
  END vss
  OBS
    LAYER met1 SPACING 0.14 ;
      RECT -2.225 0.62 769.265 9.005 ;
      RECT 766.67 -1.525 769.265 9.005 ;
      RECT 766.55 0 769.265 9.005 ;
      RECT 762.65 -1.525 765.75 9.005 ;
      RECT 760.55 0 761.85 9.005 ;
      RECT 756.65 -1.525 759.75 9.005 ;
      RECT 754.55 0 755.85 9.005 ;
      RECT 750.65 -1.525 753.75 9.005 ;
      RECT 748.55 0 749.85 9.005 ;
      RECT 744.65 -1.525 747.75 9.005 ;
      RECT 742.55 0 743.85 9.005 ;
      RECT 738.65 -1.525 741.75 9.005 ;
      RECT 736.55 0 737.85 9.005 ;
      RECT 732.65 -1.525 735.75 9.005 ;
      RECT 730.55 0 731.85 9.005 ;
      RECT 726.65 -1.525 729.75 9.005 ;
      RECT 724.55 0 725.85 9.005 ;
      RECT 720.65 -1.525 723.75 9.005 ;
      RECT 718.55 0 719.85 9.005 ;
      RECT 714.65 -1.525 717.75 9.005 ;
      RECT 712.55 0 713.85 9.005 ;
      RECT 708.65 -1.525 711.75 9.005 ;
      RECT 706.55 0 707.85 9.005 ;
      RECT 702.65 -1.525 705.75 9.005 ;
      RECT 700.55 0 701.85 9.005 ;
      RECT 696.65 -1.525 699.75 9.005 ;
      RECT 694.55 0 695.85 9.005 ;
      RECT 690.65 -1.525 693.75 9.005 ;
      RECT 688.55 0 689.85 9.005 ;
      RECT 684.65 -1.525 687.75 9.005 ;
      RECT 682.55 0 683.85 9.005 ;
      RECT 678.65 -1.525 681.75 9.005 ;
      RECT 676.55 0 677.85 9.005 ;
      RECT 672.65 -1.525 675.75 9.005 ;
      RECT 670.55 0 671.85 9.005 ;
      RECT 666.65 -1.525 669.75 9.005 ;
      RECT 664.55 0 665.85 9.005 ;
      RECT 660.65 -1.525 663.75 9.005 ;
      RECT 658.55 0 659.85 9.005 ;
      RECT 654.65 -1.525 657.75 9.005 ;
      RECT 652.55 0 653.85 9.005 ;
      RECT 648.65 -1.525 651.75 9.005 ;
      RECT 646.55 0 647.85 9.005 ;
      RECT 642.65 -1.525 645.75 9.005 ;
      RECT 640.55 0 641.85 9.005 ;
      RECT 636.65 -1.525 639.75 9.005 ;
      RECT 634.55 0 635.85 9.005 ;
      RECT 630.65 -1.525 633.75 9.005 ;
      RECT 628.55 0 629.85 9.005 ;
      RECT 624.65 -1.525 627.75 9.005 ;
      RECT 622.55 0 623.85 9.005 ;
      RECT 618.65 -1.525 621.75 9.005 ;
      RECT 616.55 0 617.85 9.005 ;
      RECT 612.65 -1.525 615.75 9.005 ;
      RECT 610.55 0 611.85 9.005 ;
      RECT 606.65 -1.525 609.75 9.005 ;
      RECT 604.55 0 605.85 9.005 ;
      RECT 600.65 -1.525 603.75 9.005 ;
      RECT 598.55 0 599.85 9.005 ;
      RECT 594.65 -1.525 597.75 9.005 ;
      RECT 592.55 0 593.85 9.005 ;
      RECT 588.65 -1.525 591.75 9.005 ;
      RECT 586.55 0 587.85 9.005 ;
      RECT 582.65 -1.525 585.75 9.005 ;
      RECT 580.55 0 581.85 9.005 ;
      RECT 576.65 -1.525 579.75 9.005 ;
      RECT 574.55 0 575.85 9.005 ;
      RECT 570.65 -1.525 573.75 9.005 ;
      RECT 568.55 0 569.85 9.005 ;
      RECT 564.65 -1.525 567.75 9.005 ;
      RECT 562.55 0 563.85 9.005 ;
      RECT 558.65 -1.525 561.75 9.005 ;
      RECT 556.55 0 557.85 9.005 ;
      RECT 552.65 -1.525 555.75 9.005 ;
      RECT 550.55 0 551.85 9.005 ;
      RECT 546.65 -1.525 549.75 9.005 ;
      RECT 544.55 0 545.85 9.005 ;
      RECT 540.65 -1.525 543.75 9.005 ;
      RECT 538.55 0 539.85 9.005 ;
      RECT 534.65 -1.525 537.75 9.005 ;
      RECT 532.55 0 533.85 9.005 ;
      RECT 528.65 -1.525 531.75 9.005 ;
      RECT 526.55 0 527.85 9.005 ;
      RECT 522.65 -1.525 525.75 9.005 ;
      RECT 520.55 0 521.85 9.005 ;
      RECT 516.65 -1.525 519.75 9.005 ;
      RECT 514.55 0 515.85 9.005 ;
      RECT 510.65 -1.525 513.75 9.005 ;
      RECT 508.55 0 509.85 9.005 ;
      RECT 504.65 -1.525 507.75 9.005 ;
      RECT 502.55 0 503.85 9.005 ;
      RECT 498.65 -1.525 501.75 9.005 ;
      RECT 496.55 0 497.85 9.005 ;
      RECT 492.65 -1.525 495.75 9.005 ;
      RECT 490.55 0 491.85 9.005 ;
      RECT 486.65 -1.525 489.75 9.005 ;
      RECT 484.55 0 485.85 9.005 ;
      RECT 480.65 -1.525 483.75 9.005 ;
      RECT 478.55 0 479.85 9.005 ;
      RECT 474.65 -1.525 477.75 9.005 ;
      RECT 472.55 0 473.85 9.005 ;
      RECT 468.65 -1.525 471.75 9.005 ;
      RECT 466.55 0 467.85 9.005 ;
      RECT 462.65 -1.525 465.75 9.005 ;
      RECT 460.55 0 461.85 9.005 ;
      RECT 456.65 -1.525 459.75 9.005 ;
      RECT 454.55 0 455.85 9.005 ;
      RECT 450.65 -1.525 453.75 9.005 ;
      RECT 448.55 0 449.85 9.005 ;
      RECT 444.65 -1.525 447.75 9.005 ;
      RECT 442.55 0 443.85 9.005 ;
      RECT 438.65 -1.525 441.75 9.005 ;
      RECT 436.55 0 437.85 9.005 ;
      RECT 432.65 -1.525 435.75 9.005 ;
      RECT 430.55 0 431.85 9.005 ;
      RECT 426.65 -1.525 429.75 9.005 ;
      RECT 424.55 0 425.85 9.005 ;
      RECT 420.65 -1.525 423.75 9.005 ;
      RECT 418.55 0 419.85 9.005 ;
      RECT 414.65 -1.525 417.75 9.005 ;
      RECT 412.55 0 413.85 9.005 ;
      RECT 408.65 -1.525 411.75 9.005 ;
      RECT 406.55 0 407.85 9.005 ;
      RECT 402.65 -1.525 405.75 9.005 ;
      RECT 400.55 0 401.85 9.005 ;
      RECT 396.65 -1.525 399.75 9.005 ;
      RECT 394.55 0 395.85 9.005 ;
      RECT 390.65 -1.525 393.75 9.005 ;
      RECT 388.55 0 389.85 9.005 ;
      RECT 384.65 -1.525 387.75 9.005 ;
      RECT 382.55 0 383.85 9.005 ;
      RECT 378.65 -1.525 381.75 9.005 ;
      RECT 376.55 0 377.85 9.005 ;
      RECT 372.65 -1.525 375.75 9.005 ;
      RECT 370.55 0 371.85 9.005 ;
      RECT 366.65 -1.525 369.75 9.005 ;
      RECT 364.55 0 365.85 9.005 ;
      RECT 360.65 -1.525 363.75 9.005 ;
      RECT 358.55 0 359.85 9.005 ;
      RECT 354.65 -1.525 357.75 9.005 ;
      RECT 352.55 0 353.85 9.005 ;
      RECT 348.65 -1.525 351.75 9.005 ;
      RECT 346.55 0 347.85 9.005 ;
      RECT 342.65 -1.525 345.75 9.005 ;
      RECT 340.55 0 341.85 9.005 ;
      RECT 336.65 -1.525 339.75 9.005 ;
      RECT 334.55 0 335.85 9.005 ;
      RECT 330.65 -1.525 333.75 9.005 ;
      RECT 328.55 0 329.85 9.005 ;
      RECT 324.65 -1.525 327.75 9.005 ;
      RECT 322.55 0 323.85 9.005 ;
      RECT 318.65 -1.525 321.75 9.005 ;
      RECT 316.55 0 317.85 9.005 ;
      RECT 312.65 -1.525 315.75 9.005 ;
      RECT 310.55 0 311.85 9.005 ;
      RECT 306.65 -1.525 309.75 9.005 ;
      RECT 304.55 0 305.85 9.005 ;
      RECT 300.65 -1.525 303.75 9.005 ;
      RECT 298.55 0 299.85 9.005 ;
      RECT 294.65 -1.525 297.75 9.005 ;
      RECT 292.55 0 293.85 9.005 ;
      RECT 288.65 -1.525 291.75 9.005 ;
      RECT 286.55 0 287.85 9.005 ;
      RECT 282.65 -1.525 285.75 9.005 ;
      RECT 280.55 0 281.85 9.005 ;
      RECT 276.65 -1.525 279.75 9.005 ;
      RECT 274.55 0 275.85 9.005 ;
      RECT 270.65 -1.525 273.75 9.005 ;
      RECT 268.55 0 269.85 9.005 ;
      RECT 264.65 -1.525 267.75 9.005 ;
      RECT 262.55 0 263.85 9.005 ;
      RECT 258.65 -1.525 261.75 9.005 ;
      RECT 256.55 0 257.85 9.005 ;
      RECT 252.65 -1.525 255.75 9.005 ;
      RECT 250.55 0 251.85 9.005 ;
      RECT 246.65 -1.525 249.75 9.005 ;
      RECT 244.55 0 245.85 9.005 ;
      RECT 240.65 -1.525 243.75 9.005 ;
      RECT 238.55 0 239.85 9.005 ;
      RECT 234.65 -1.525 237.75 9.005 ;
      RECT 232.55 0 233.85 9.005 ;
      RECT 228.65 -1.525 231.75 9.005 ;
      RECT 226.55 0 227.85 9.005 ;
      RECT 222.65 -1.525 225.75 9.005 ;
      RECT 220.55 0 221.85 9.005 ;
      RECT 216.65 -1.525 219.75 9.005 ;
      RECT 214.55 0 215.85 9.005 ;
      RECT 210.65 -1.525 213.75 9.005 ;
      RECT 208.55 0 209.85 9.005 ;
      RECT 204.65 -1.525 207.75 9.005 ;
      RECT 202.55 0 203.85 9.005 ;
      RECT 198.65 -1.525 201.75 9.005 ;
      RECT 196.55 0 197.85 9.005 ;
      RECT 192.65 -1.525 195.75 9.005 ;
      RECT 190.55 0 191.85 9.005 ;
      RECT 186.65 -1.525 189.75 9.005 ;
      RECT 184.55 0 185.85 9.005 ;
      RECT 180.65 -1.525 183.75 9.005 ;
      RECT 178.55 0 179.85 9.005 ;
      RECT 174.65 -1.525 177.75 9.005 ;
      RECT 172.55 0 173.85 9.005 ;
      RECT 168.65 -1.525 171.75 9.005 ;
      RECT 166.55 0 167.85 9.005 ;
      RECT 162.65 -1.525 165.75 9.005 ;
      RECT 160.55 0 161.85 9.005 ;
      RECT 156.65 -1.525 159.75 9.005 ;
      RECT 154.55 0 155.85 9.005 ;
      RECT 150.65 -1.525 153.75 9.005 ;
      RECT 148.55 0 149.85 9.005 ;
      RECT 144.65 -1.525 147.75 9.005 ;
      RECT 142.55 0 143.85 9.005 ;
      RECT 138.65 -1.525 141.75 9.005 ;
      RECT 136.55 0 137.85 9.005 ;
      RECT 132.65 -1.525 135.75 9.005 ;
      RECT 130.55 0 131.85 9.005 ;
      RECT 126.65 -1.525 129.75 9.005 ;
      RECT 124.55 0 125.85 9.005 ;
      RECT 120.65 -1.525 123.75 9.005 ;
      RECT 118.55 0 119.85 9.005 ;
      RECT 114.65 -1.525 117.75 9.005 ;
      RECT 112.55 0 113.85 9.005 ;
      RECT 108.65 -1.525 111.75 9.005 ;
      RECT 106.55 0 107.85 9.005 ;
      RECT 102.65 -1.525 105.75 9.005 ;
      RECT 100.55 0 101.85 9.005 ;
      RECT 96.65 -1.525 99.75 9.005 ;
      RECT 94.55 0 95.85 9.005 ;
      RECT 90.65 -1.525 93.75 9.005 ;
      RECT 88.55 0 89.85 9.005 ;
      RECT 84.65 -1.525 87.75 9.005 ;
      RECT 82.55 0 83.85 9.005 ;
      RECT 78.65 -1.525 81.75 9.005 ;
      RECT 76.55 0 77.85 9.005 ;
      RECT 72.65 -1.525 75.75 9.005 ;
      RECT 70.55 0 71.85 9.005 ;
      RECT 66.65 -1.525 69.75 9.005 ;
      RECT 64.55 0 65.85 9.005 ;
      RECT 60.65 -1.525 63.75 9.005 ;
      RECT 58.55 0 59.85 9.005 ;
      RECT 54.65 -1.525 57.75 9.005 ;
      RECT 52.55 0 53.85 9.005 ;
      RECT 48.65 -1.525 51.75 9.005 ;
      RECT 46.55 0 47.85 9.005 ;
      RECT 42.65 -1.525 45.75 9.005 ;
      RECT 40.55 0 41.85 9.005 ;
      RECT 36.65 -1.525 39.75 9.005 ;
      RECT 34.55 0 35.85 9.005 ;
      RECT 30.65 -1.525 33.75 9.005 ;
      RECT 28.55 0 29.85 9.005 ;
      RECT 24.65 -1.525 27.75 9.005 ;
      RECT 22.55 0 23.85 9.005 ;
      RECT 18.65 -1.525 21.75 9.005 ;
      RECT 16.55 0 17.85 9.005 ;
      RECT 12.65 -1.525 15.75 9.005 ;
      RECT 10.55 0 11.85 9.005 ;
      RECT 6.65 -1.525 9.75 9.005 ;
      RECT 4.67 0 5.85 9.005 ;
      RECT 2.14 -1.525 3.75 9.005 ;
      RECT 0.65 -1.525 1.22 9.005 ;
      RECT -2.225 -1.525 -0.77 9.005 ;
      RECT 760.67 -1.525 761.73 9.005 ;
      RECT 754.67 -1.525 755.73 9.005 ;
      RECT 748.67 -1.525 749.73 9.005 ;
      RECT 742.67 -1.525 743.73 9.005 ;
      RECT 736.67 -1.525 737.73 9.005 ;
      RECT 730.67 -1.525 731.73 9.005 ;
      RECT 724.67 -1.525 725.73 9.005 ;
      RECT 718.67 -1.525 719.73 9.005 ;
      RECT 712.67 -1.525 713.73 9.005 ;
      RECT 706.67 -1.525 707.73 9.005 ;
      RECT 700.67 -1.525 701.73 9.005 ;
      RECT 694.67 -1.525 695.73 9.005 ;
      RECT 688.67 -1.525 689.73 9.005 ;
      RECT 682.67 -1.525 683.73 9.005 ;
      RECT 676.67 -1.525 677.73 9.005 ;
      RECT 670.67 -1.525 671.73 9.005 ;
      RECT 664.67 -1.525 665.73 9.005 ;
      RECT 658.67 -1.525 659.73 9.005 ;
      RECT 652.67 -1.525 653.73 9.005 ;
      RECT 646.67 -1.525 647.73 9.005 ;
      RECT 640.67 -1.525 641.73 9.005 ;
      RECT 634.67 -1.525 635.73 9.005 ;
      RECT 628.67 -1.525 629.73 9.005 ;
      RECT 622.67 -1.525 623.73 9.005 ;
      RECT 616.67 -1.525 617.73 9.005 ;
      RECT 610.67 -1.525 611.73 9.005 ;
      RECT 604.67 -1.525 605.73 9.005 ;
      RECT 598.67 -1.525 599.73 9.005 ;
      RECT 592.67 -1.525 593.73 9.005 ;
      RECT 586.67 -1.525 587.73 9.005 ;
      RECT 580.67 -1.525 581.73 9.005 ;
      RECT 574.67 -1.525 575.73 9.005 ;
      RECT 568.67 -1.525 569.73 9.005 ;
      RECT 562.67 -1.525 563.73 9.005 ;
      RECT 556.67 -1.525 557.73 9.005 ;
      RECT 550.67 -1.525 551.73 9.005 ;
      RECT 544.67 -1.525 545.73 9.005 ;
      RECT 538.67 -1.525 539.73 9.005 ;
      RECT 532.67 -1.525 533.73 9.005 ;
      RECT 526.67 -1.525 527.73 9.005 ;
      RECT 520.67 -1.525 521.73 9.005 ;
      RECT 514.67 -1.525 515.73 9.005 ;
      RECT 508.67 -1.525 509.73 9.005 ;
      RECT 502.67 -1.525 503.73 9.005 ;
      RECT 496.67 -1.525 497.73 9.005 ;
      RECT 490.67 -1.525 491.73 9.005 ;
      RECT 484.67 -1.525 485.73 9.005 ;
      RECT 478.67 -1.525 479.73 9.005 ;
      RECT 472.67 -1.525 473.73 9.005 ;
      RECT 466.67 -1.525 467.73 9.005 ;
      RECT 460.67 -1.525 461.73 9.005 ;
      RECT 454.67 -1.525 455.73 9.005 ;
      RECT 448.67 -1.525 449.73 9.005 ;
      RECT 442.67 -1.525 443.73 9.005 ;
      RECT 436.67 -1.525 437.73 9.005 ;
      RECT 430.67 -1.525 431.73 9.005 ;
      RECT 424.67 -1.525 425.73 9.005 ;
      RECT 418.67 -1.525 419.73 9.005 ;
      RECT 412.67 -1.525 413.73 9.005 ;
      RECT 406.67 -1.525 407.73 9.005 ;
      RECT 400.67 -1.525 401.73 9.005 ;
      RECT 394.67 -1.525 395.73 9.005 ;
      RECT 388.67 -1.525 389.73 9.005 ;
      RECT 382.67 -1.525 383.73 9.005 ;
      RECT 376.67 -1.525 377.73 9.005 ;
      RECT 370.67 -1.525 371.73 9.005 ;
      RECT 364.67 -1.525 365.73 9.005 ;
      RECT 358.67 -1.525 359.73 9.005 ;
      RECT 352.67 -1.525 353.73 9.005 ;
      RECT 346.67 -1.525 347.73 9.005 ;
      RECT 340.67 -1.525 341.73 9.005 ;
      RECT 334.67 -1.525 335.73 9.005 ;
      RECT 328.67 -1.525 329.73 9.005 ;
      RECT 322.67 -1.525 323.73 9.005 ;
      RECT 316.67 -1.525 317.73 9.005 ;
      RECT 310.67 -1.525 311.73 9.005 ;
      RECT 304.67 -1.525 305.73 9.005 ;
      RECT 298.67 -1.525 299.73 9.005 ;
      RECT 292.67 -1.525 293.73 9.005 ;
      RECT 286.67 -1.525 287.73 9.005 ;
      RECT 280.67 -1.525 281.73 9.005 ;
      RECT 274.67 -1.525 275.73 9.005 ;
      RECT 268.67 -1.525 269.73 9.005 ;
      RECT 262.67 -1.525 263.73 9.005 ;
      RECT 256.67 -1.525 257.73 9.005 ;
      RECT 250.67 -1.525 251.73 9.005 ;
      RECT 244.67 -1.525 245.73 9.005 ;
      RECT 238.67 -1.525 239.73 9.005 ;
      RECT 232.67 -1.525 233.73 9.005 ;
      RECT 226.67 -1.525 227.73 9.005 ;
      RECT 220.67 -1.525 221.73 9.005 ;
      RECT 214.67 -1.525 215.73 9.005 ;
      RECT 208.67 -1.525 209.73 9.005 ;
      RECT 202.67 -1.525 203.73 9.005 ;
      RECT 196.67 -1.525 197.73 9.005 ;
      RECT 190.67 -1.525 191.73 9.005 ;
      RECT 184.67 -1.525 185.73 9.005 ;
      RECT 178.67 -1.525 179.73 9.005 ;
      RECT 172.67 -1.525 173.73 9.005 ;
      RECT 166.67 -1.525 167.73 9.005 ;
      RECT 160.67 -1.525 161.73 9.005 ;
      RECT 154.67 -1.525 155.73 9.005 ;
      RECT 148.67 -1.525 149.73 9.005 ;
      RECT 142.67 -1.525 143.73 9.005 ;
      RECT 136.67 -1.525 137.73 9.005 ;
      RECT 130.67 -1.525 131.73 9.005 ;
      RECT 124.67 -1.525 125.73 9.005 ;
      RECT 118.67 -1.525 119.73 9.005 ;
      RECT 112.67 -1.525 113.73 9.005 ;
      RECT 106.67 -1.525 107.73 9.005 ;
      RECT 100.67 -1.525 101.73 9.005 ;
      RECT 94.67 -1.525 95.73 9.005 ;
      RECT 88.67 -1.525 89.73 9.005 ;
      RECT 82.67 -1.525 83.73 9.005 ;
      RECT 76.67 -1.525 77.73 9.005 ;
      RECT 70.67 -1.525 71.73 9.005 ;
      RECT 64.67 -1.525 65.73 9.005 ;
      RECT 58.67 -1.525 59.73 9.005 ;
      RECT 52.67 -1.525 53.73 9.005 ;
      RECT 46.67 -1.525 47.73 9.005 ;
      RECT 40.67 -1.525 41.73 9.005 ;
      RECT 34.67 -1.525 35.73 9.005 ;
      RECT 28.67 -1.525 29.73 9.005 ;
      RECT 22.67 -1.525 23.73 9.005 ;
      RECT 16.67 -1.525 17.73 9.005 ;
      RECT 10.67 -1.525 11.73 9.005 ;
      RECT 4.67 -1.525 5.73 9.005 ;
      RECT -2.225 -1.525 769.265 -0.3 ;
    LAYER met2 ;
      RECT -2.2 -1.52 769.24 -1.2 ;
      RECT -2.225 -1.5 769.265 -1.22 ;
      RECT -2.2 -0.16 769.24 0.16 ;
      RECT -2.225 -0.14 769.265 0.14 ;
      RECT -2.2 1.2 769.24 1.52 ;
      RECT -2.225 1.22 769.265 1.5 ;
      RECT -2.2 2.56 769.24 2.88 ;
      RECT -2.225 2.58 769.265 2.86 ;
      RECT 764.84 3.92 769.24 4.24 ;
      RECT 764.84 3.94 769.265 4.22 ;
      RECT 762.8 5.28 769.24 5.6 ;
      RECT 762.8 5.3 769.265 5.58 ;
      RECT 767.56 6.64 769.24 6.96 ;
      RECT 767.56 6.66 769.265 6.94 ;
      RECT -2.2 8 769.24 8.32 ;
      RECT -2.225 8.02 769.265 8.3 ;
      RECT -2.2 5.28 3.56 5.6 ;
      RECT -2.225 5.3 3.56 5.58 ;
      RECT -2.2 3.92 0.84 4.24 ;
      RECT -2.225 3.94 0.84 4.22 ;
      RECT -2.2 6.64 -0.52 6.96 ;
      RECT -2.225 6.66 -0.52 6.94 ;
      RECT -2.2 -0.84 769.24 -0.52 ;
      RECT -2.2 0.52 769.24 0.84 ;
      RECT -2.2 1.88 769.24 2.2 ;
      RECT 759.4 3.24 769.24 3.56 ;
      RECT 764.84 4.6 769.24 4.92 ;
      RECT 767.56 5.96 769.24 6.28 ;
      RECT -2.2 7.32 769.24 7.64 ;
      RECT -2.2 8.68 769.24 9 ;
      RECT -2.2 3.24 6.96 3.56 ;
      RECT -2.2 4.6 0.84 4.92 ;
      RECT -2.2 5.96 -0.52 6.28 ;
    LAYER met2 SPACING 0.14 ;
      RECT -2.225 0.52 769.265 9.005 ;
      RECT 766.67 -1.525 769.265 9.005 ;
      RECT 762.65 -1.525 765.75 9.005 ;
      RECT 760.67 -1.525 761.73 9.005 ;
      RECT 756.65 -1.525 759.75 9.005 ;
      RECT 754.67 -1.525 755.73 9.005 ;
      RECT 750.65 -1.525 753.75 9.005 ;
      RECT 748.67 -1.525 749.73 9.005 ;
      RECT 744.65 -1.525 747.75 9.005 ;
      RECT 742.67 -1.525 743.73 9.005 ;
      RECT 738.65 -1.525 741.75 9.005 ;
      RECT 736.67 -1.525 737.73 9.005 ;
      RECT 732.65 -1.525 735.75 9.005 ;
      RECT 730.67 -1.525 731.73 9.005 ;
      RECT 726.65 -1.525 729.75 9.005 ;
      RECT 724.67 -1.525 725.73 9.005 ;
      RECT 720.65 -1.525 723.75 9.005 ;
      RECT 718.67 -1.525 719.73 9.005 ;
      RECT 714.65 -1.525 717.75 9.005 ;
      RECT 712.67 -1.525 713.73 9.005 ;
      RECT 708.65 -1.525 711.75 9.005 ;
      RECT 706.67 -1.525 707.73 9.005 ;
      RECT 702.65 -1.525 705.75 9.005 ;
      RECT 700.67 -1.525 701.73 9.005 ;
      RECT 696.65 -1.525 699.75 9.005 ;
      RECT 694.67 -1.525 695.73 9.005 ;
      RECT 690.65 -1.525 693.75 9.005 ;
      RECT 688.67 -1.525 689.73 9.005 ;
      RECT 684.65 -1.525 687.75 9.005 ;
      RECT 682.67 -1.525 683.73 9.005 ;
      RECT 678.65 -1.525 681.75 9.005 ;
      RECT 676.67 -1.525 677.73 9.005 ;
      RECT 672.65 -1.525 675.75 9.005 ;
      RECT 670.67 -1.525 671.73 9.005 ;
      RECT 666.65 -1.525 669.75 9.005 ;
      RECT 664.67 -1.525 665.73 9.005 ;
      RECT 660.65 -1.525 663.75 9.005 ;
      RECT 658.67 -1.525 659.73 9.005 ;
      RECT 654.65 -1.525 657.75 9.005 ;
      RECT 652.67 -1.525 653.73 9.005 ;
      RECT 648.65 -1.525 651.75 9.005 ;
      RECT 646.67 -1.525 647.73 9.005 ;
      RECT 642.65 -1.525 645.75 9.005 ;
      RECT 640.67 -1.525 641.73 9.005 ;
      RECT 636.65 -1.525 639.75 9.005 ;
      RECT 634.67 -1.525 635.73 9.005 ;
      RECT 630.65 -1.525 633.75 9.005 ;
      RECT 628.67 -1.525 629.73 9.005 ;
      RECT 624.65 -1.525 627.75 9.005 ;
      RECT 622.67 -1.525 623.73 9.005 ;
      RECT 618.65 -1.525 621.75 9.005 ;
      RECT 616.67 -1.525 617.73 9.005 ;
      RECT 612.65 -1.525 615.75 9.005 ;
      RECT 610.67 -1.525 611.73 9.005 ;
      RECT 606.65 -1.525 609.75 9.005 ;
      RECT 604.67 -1.525 605.73 9.005 ;
      RECT 600.65 -1.525 603.75 9.005 ;
      RECT 598.67 -1.525 599.73 9.005 ;
      RECT 594.65 -1.525 597.75 9.005 ;
      RECT 592.67 -1.525 593.73 9.005 ;
      RECT 588.65 -1.525 591.75 9.005 ;
      RECT 586.67 -1.525 587.73 9.005 ;
      RECT 582.65 -1.525 585.75 9.005 ;
      RECT 580.67 -1.525 581.73 9.005 ;
      RECT 576.65 -1.525 579.75 9.005 ;
      RECT 574.67 -1.525 575.73 9.005 ;
      RECT 570.65 -1.525 573.75 9.005 ;
      RECT 568.67 -1.525 569.73 9.005 ;
      RECT 564.65 -1.525 567.75 9.005 ;
      RECT 562.67 -1.525 563.73 9.005 ;
      RECT 558.65 -1.525 561.75 9.005 ;
      RECT 556.67 -1.525 557.73 9.005 ;
      RECT 552.65 -1.525 555.75 9.005 ;
      RECT 550.67 -1.525 551.73 9.005 ;
      RECT 546.65 -1.525 549.75 9.005 ;
      RECT 544.67 -1.525 545.73 9.005 ;
      RECT 540.65 -1.525 543.75 9.005 ;
      RECT 538.67 -1.525 539.73 9.005 ;
      RECT 534.65 -1.525 537.75 9.005 ;
      RECT 532.67 -1.525 533.73 9.005 ;
      RECT 528.65 -1.525 531.75 9.005 ;
      RECT 526.67 -1.525 527.73 9.005 ;
      RECT 522.65 -1.525 525.75 9.005 ;
      RECT 520.67 -1.525 521.73 9.005 ;
      RECT 516.65 -1.525 519.75 9.005 ;
      RECT 514.67 -1.525 515.73 9.005 ;
      RECT 510.65 -1.525 513.75 9.005 ;
      RECT 508.67 -1.525 509.73 9.005 ;
      RECT 504.65 -1.525 507.75 9.005 ;
      RECT 502.67 -1.525 503.73 9.005 ;
      RECT 498.65 -1.525 501.75 9.005 ;
      RECT 496.67 -1.525 497.73 9.005 ;
      RECT 492.65 -1.525 495.75 9.005 ;
      RECT 490.67 -1.525 491.73 9.005 ;
      RECT 486.65 -1.525 489.75 9.005 ;
      RECT 484.67 -1.525 485.73 9.005 ;
      RECT 480.65 -1.525 483.75 9.005 ;
      RECT 478.67 -1.525 479.73 9.005 ;
      RECT 474.65 -1.525 477.75 9.005 ;
      RECT 472.67 -1.525 473.73 9.005 ;
      RECT 468.65 -1.525 471.75 9.005 ;
      RECT 466.67 -1.525 467.73 9.005 ;
      RECT 462.65 -1.525 465.75 9.005 ;
      RECT 460.67 -1.525 461.73 9.005 ;
      RECT 456.65 -1.525 459.75 9.005 ;
      RECT 454.67 -1.525 455.73 9.005 ;
      RECT 450.65 -1.525 453.75 9.005 ;
      RECT 448.67 -1.525 449.73 9.005 ;
      RECT 444.65 -1.525 447.75 9.005 ;
      RECT 442.67 -1.525 443.73 9.005 ;
      RECT 438.65 -1.525 441.75 9.005 ;
      RECT 436.67 -1.525 437.73 9.005 ;
      RECT 432.65 -1.525 435.75 9.005 ;
      RECT 430.67 -1.525 431.73 9.005 ;
      RECT 426.65 -1.525 429.75 9.005 ;
      RECT 424.67 -1.525 425.73 9.005 ;
      RECT 420.65 -1.525 423.75 9.005 ;
      RECT 418.67 -1.525 419.73 9.005 ;
      RECT 414.65 -1.525 417.75 9.005 ;
      RECT 412.67 -1.525 413.73 9.005 ;
      RECT 408.65 -1.525 411.75 9.005 ;
      RECT 406.67 -1.525 407.73 9.005 ;
      RECT 402.65 -1.525 405.75 9.005 ;
      RECT 400.67 -1.525 401.73 9.005 ;
      RECT 396.65 -1.525 399.75 9.005 ;
      RECT 394.67 -1.525 395.73 9.005 ;
      RECT 390.65 -1.525 393.75 9.005 ;
      RECT 388.67 -1.525 389.73 9.005 ;
      RECT 384.65 -1.525 387.75 9.005 ;
      RECT 382.67 -1.525 383.73 9.005 ;
      RECT 378.65 -1.525 381.75 9.005 ;
      RECT 376.67 -1.525 377.73 9.005 ;
      RECT 372.65 -1.525 375.75 9.005 ;
      RECT 370.67 -1.525 371.73 9.005 ;
      RECT 366.65 -1.525 369.75 9.005 ;
      RECT 364.67 -1.525 365.73 9.005 ;
      RECT 360.65 -1.525 363.75 9.005 ;
      RECT 358.67 -1.525 359.73 9.005 ;
      RECT 354.65 -1.525 357.75 9.005 ;
      RECT 352.67 -1.525 353.73 9.005 ;
      RECT 348.65 -1.525 351.75 9.005 ;
      RECT 346.67 -1.525 347.73 9.005 ;
      RECT 342.65 -1.525 345.75 9.005 ;
      RECT 340.67 -1.525 341.73 9.005 ;
      RECT 336.65 -1.525 339.75 9.005 ;
      RECT 334.67 -1.525 335.73 9.005 ;
      RECT 330.65 -1.525 333.75 9.005 ;
      RECT 328.67 -1.525 329.73 9.005 ;
      RECT 324.65 -1.525 327.75 9.005 ;
      RECT 322.67 -1.525 323.73 9.005 ;
      RECT 318.65 -1.525 321.75 9.005 ;
      RECT 316.67 -1.525 317.73 9.005 ;
      RECT 312.65 -1.525 315.75 9.005 ;
      RECT 310.67 -1.525 311.73 9.005 ;
      RECT 306.65 -1.525 309.75 9.005 ;
      RECT 304.67 -1.525 305.73 9.005 ;
      RECT 300.65 -1.525 303.75 9.005 ;
      RECT 298.67 -1.525 299.73 9.005 ;
      RECT 294.65 -1.525 297.75 9.005 ;
      RECT 292.67 -1.525 293.73 9.005 ;
      RECT 288.65 -1.525 291.75 9.005 ;
      RECT 286.67 -1.525 287.73 9.005 ;
      RECT 282.65 -1.525 285.75 9.005 ;
      RECT 280.67 -1.525 281.73 9.005 ;
      RECT 276.65 -1.525 279.75 9.005 ;
      RECT 274.67 -1.525 275.73 9.005 ;
      RECT 270.65 -1.525 273.75 9.005 ;
      RECT 268.67 -1.525 269.73 9.005 ;
      RECT 264.65 -1.525 267.75 9.005 ;
      RECT 262.67 -1.525 263.73 9.005 ;
      RECT 258.65 -1.525 261.75 9.005 ;
      RECT 256.67 -1.525 257.73 9.005 ;
      RECT 252.65 -1.525 255.75 9.005 ;
      RECT 250.67 -1.525 251.73 9.005 ;
      RECT 246.65 -1.525 249.75 9.005 ;
      RECT 244.67 -1.525 245.73 9.005 ;
      RECT 240.65 -1.525 243.75 9.005 ;
      RECT 238.67 -1.525 239.73 9.005 ;
      RECT 234.65 -1.525 237.75 9.005 ;
      RECT 232.67 -1.525 233.73 9.005 ;
      RECT 228.65 -1.525 231.75 9.005 ;
      RECT 226.67 -1.525 227.73 9.005 ;
      RECT 222.65 -1.525 225.75 9.005 ;
      RECT 220.67 -1.525 221.73 9.005 ;
      RECT 216.65 -1.525 219.75 9.005 ;
      RECT 214.67 -1.525 215.73 9.005 ;
      RECT 210.65 -1.525 213.75 9.005 ;
      RECT 208.67 -1.525 209.73 9.005 ;
      RECT 204.65 -1.525 207.75 9.005 ;
      RECT 202.67 -1.525 203.73 9.005 ;
      RECT 198.65 -1.525 201.75 9.005 ;
      RECT 196.67 -1.525 197.73 9.005 ;
      RECT 192.65 -1.525 195.75 9.005 ;
      RECT 190.67 -1.525 191.73 9.005 ;
      RECT 186.65 -1.525 189.75 9.005 ;
      RECT 184.67 -1.525 185.73 9.005 ;
      RECT 180.65 -1.525 183.75 9.005 ;
      RECT 178.67 -1.525 179.73 9.005 ;
      RECT 174.65 -1.525 177.75 9.005 ;
      RECT 172.67 -1.525 173.73 9.005 ;
      RECT 168.65 -1.525 171.75 9.005 ;
      RECT 166.67 -1.525 167.73 9.005 ;
      RECT 162.65 -1.525 165.75 9.005 ;
      RECT 160.67 -1.525 161.73 9.005 ;
      RECT 156.65 -1.525 159.75 9.005 ;
      RECT 154.67 -1.525 155.73 9.005 ;
      RECT 150.65 -1.525 153.75 9.005 ;
      RECT 148.67 -1.525 149.73 9.005 ;
      RECT 144.65 -1.525 147.75 9.005 ;
      RECT 142.67 -1.525 143.73 9.005 ;
      RECT 138.65 -1.525 141.75 9.005 ;
      RECT 136.67 -1.525 137.73 9.005 ;
      RECT 132.65 -1.525 135.75 9.005 ;
      RECT 130.67 -1.525 131.73 9.005 ;
      RECT 126.65 -1.525 129.75 9.005 ;
      RECT 124.67 -1.525 125.73 9.005 ;
      RECT 120.65 -1.525 123.75 9.005 ;
      RECT 118.67 -1.525 119.73 9.005 ;
      RECT 114.65 -1.525 117.75 9.005 ;
      RECT 112.67 -1.525 113.73 9.005 ;
      RECT 108.65 -1.525 111.75 9.005 ;
      RECT 106.67 -1.525 107.73 9.005 ;
      RECT 102.65 -1.525 105.75 9.005 ;
      RECT 100.67 -1.525 101.73 9.005 ;
      RECT 96.65 -1.525 99.75 9.005 ;
      RECT 94.67 -1.525 95.73 9.005 ;
      RECT 90.65 -1.525 93.75 9.005 ;
      RECT 88.67 -1.525 89.73 9.005 ;
      RECT 84.65 -1.525 87.75 9.005 ;
      RECT 82.67 -1.525 83.73 9.005 ;
      RECT 78.65 -1.525 81.75 9.005 ;
      RECT 76.67 -1.525 77.73 9.005 ;
      RECT 72.65 -1.525 75.75 9.005 ;
      RECT 70.67 -1.525 71.73 9.005 ;
      RECT 66.65 -1.525 69.75 9.005 ;
      RECT 64.67 -1.525 65.73 9.005 ;
      RECT 60.65 -1.525 63.75 9.005 ;
      RECT 58.67 -1.525 59.73 9.005 ;
      RECT 54.65 -1.525 57.75 9.005 ;
      RECT 52.67 -1.525 53.73 9.005 ;
      RECT 48.65 -1.525 51.75 9.005 ;
      RECT 46.67 -1.525 47.73 9.005 ;
      RECT 42.65 -1.525 45.75 9.005 ;
      RECT 40.67 -1.525 41.73 9.005 ;
      RECT 36.65 -1.525 39.75 9.005 ;
      RECT 34.67 -1.525 35.73 9.005 ;
      RECT 30.65 -1.525 33.75 9.005 ;
      RECT 28.67 -1.525 29.73 9.005 ;
      RECT 24.65 -1.525 27.75 9.005 ;
      RECT 22.67 -1.525 23.73 9.005 ;
      RECT 18.65 -1.525 21.75 9.005 ;
      RECT 16.67 -1.525 17.73 9.005 ;
      RECT 12.65 -1.525 15.75 9.005 ;
      RECT 10.67 -1.525 11.73 9.005 ;
      RECT 6.65 -1.525 9.75 9.005 ;
      RECT 4.67 -1.525 5.73 9.005 ;
      RECT 2.14 -1.525 3.75 9.005 ;
      RECT 0.65 -1.525 1.22 9.005 ;
      RECT -2.225 -1.525 -0.77 9.005 ;
      RECT -2.225 -1.525 769.265 0.16 ;
  END
END tristate_inv_delay_line_128

END LIBRARY
